/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */
/* With case-insensitive names (SPICE-compatible) */

module spm(
    inout vpwr,
    inout vgnd,
    input clk,
    output p,
    input rst,
    input y,
    input VDD,
    input VSS,
    input [31:0] x
);

wire p ;
wire [31:0] x ;
wire y ;
wire _168_ ;
wire \pp[29]  ;
wire _321_ ;
wire _130_ ;
wire _224_ ;
wire _033_ ;
wire _262_ ;
wire _318_ ;
wire _071_ ;
wire _127_ ;
wire _165_ ;
wire _259_ ;
wire _068_ ;
wire _297_ ;
wire \pp[19]  ;
wire _221_ ;
wire _030_ ;
wire _315_ ;
wire \pp[6]  ;
wire _124_ ;
wire _162_ ;
wire _218_ ;
wire _027_ ;
wire _256_ ;
wire _065_ ;
wire _294_ ;
wire _159_ ;
wire _197_ ;
wire _312_ ;
wire _121_ ;
wire clk_0_48 ;
wire _215_ ;
wire _024_ ;
wire _253_ ;
wire _309_ ;
wire _062_ ;
wire _118_ ;
wire _291_ ;
wire _156_ ;
wire \pp[24]  ;
wire _194_ ;
wire _059_ ;
wire _288_ ;
wire _097_ ;
wire clk_0_16 ;
wire _212_ ;
wire _021_ ;
wire _250_ ;
wire _306_ ;
wire _115_ ;
wire _153_ ;
wire _209_ ;
wire _018_ ;
wire _191_ ;
wire _247_ ;
wire _056_ ;
wire \pp[14]  ;
wire _285_ ;
wire _094_ ;
wire _188_ ;
wire \tcmp.s  ;
wire _303_ ;
wire _112_ ;
wire clk ;
wire _150_ ;
wire _206_ ;
wire _015_ ;
wire _244_ ;
wire _053_ ;
wire _109_ ;
wire _282_ ;
wire _091_ ;
wire _147_ ;
wire _185_ ;
wire \csa0.sc  ;
wire _279_ ;
wire _088_ ;
wire _300_ ;
wire _203_ ;
wire _012_ ;
wire _241_ ;
wire _050_ ;
wire _106_ ;
wire \pp[8]  ;
wire _144_ ;
wire _009_ ;
wire _182_ ;
wire _238_ ;
wire _047_ ;
wire _276_ ;
wire _085_ ;
wire _179_ ;
wire _200_ ;
wire VSS ;
wire _103_ ;
wire _141_ ;
wire _006_ ;
wire _235_ ;
wire _044_ ;
wire _273_ ;
wire _329_ ;
wire _082_ ;
wire _138_ ;
wire _176_ ;
wire \pp[26]  ;
wire _079_ ;
wire _100_ ;
wire _003_ ;
wire _232_ ;
wire _041_ ;
wire _270_ ;
wire _326_ ;
wire _135_ ;
wire _173_ ;
wire _229_ ;
wire _038_ ;
wire _267_ ;
wire _076_ ;
wire \csa0.hsum2  ;
wire \pp[16]  ;
wire _000_ ;
wire \pp[3]  ;
wire _323_ ;
wire _132_ ;
wire _170_ ;
wire _226_ ;
wire _035_ ;
wire _264_ ;
wire _073_ ;
wire _129_ ;
wire _167_ ;
wire _299_ ;
wire _320_ ;
wire _223_ ;
wire _032_ ;
wire _261_ ;
wire _317_ ;
wire _070_ ;
wire _126_ ;
wire \pp[21]  ;
wire _164_ ;
wire _029_ ;
wire _258_ ;
wire _067_ ;
wire _296_ ;
wire clk_0_0 ;
wire _199_ ;
wire _220_ ;
wire _314_ ;
wire VDD ;
wire _123_ ;
wire _161_ ;
wire _217_ ;
wire _026_ ;
wire \pp[11]  ;
wire _255_ ;
wire _064_ ;
wire _293_ ;
wire _158_ ;
wire _196_ ;
wire \pp[28]  ;
wire _099_ ;
wire _311_ ;
wire _120_ ;
wire clk_0_32 ;
wire _214_ ;
wire _023_ ;
wire _252_ ;
wire _308_ ;
wire _061_ ;
wire _117_ ;
wire rst ;
wire _290_ ;
wire _155_ ;
wire _193_ ;
wire _249_ ;
wire _058_ ;
wire _287_ ;
wire _096_ ;
wire \pp[18]  ;
wire _211_ ;
wire _020_ ;
wire _305_ ;
wire \pp[5]  ;
wire _114_ ;
wire _152_ ;
wire _208_ ;
wire _017_ ;
wire _190_ ;
wire _246_ ;
wire _055_ ;
wire _284_ ;
wire _093_ ;
wire _149_ ;
wire _187_ ;
wire _302_ ;
wire _111_ ;
wire _205_ ;
wire _014_ ;
wire _243_ ;
wire _052_ ;
wire _108_ ;
wire _281_ ;
wire _090_ ;
wire _146_ ;
wire \pp[23]  ;
wire _184_ ;
wire _049_ ;
wire _278_ ;
wire _087_ ;
wire _202_ ;
wire _011_ ;
wire _240_ ;
wire _105_ ;
wire _143_ ;
wire _008_ ;
wire _181_ ;
wire _237_ ;
wire _046_ ;
wire \pp[13]  ;
wire _275_ ;
wire _084_ ;
wire _178_ ;
wire _102_ ;
wire _140_ ;
wire _005_ ;
wire _234_ ;
wire _043_ ;
wire _272_ ;
wire _328_ ;
wire _081_ ;
wire _137_ ;
wire _175_ ;
wire _269_ ;
wire _078_ ;
wire _002_ ;
wire _231_ ;
wire _040_ ;
wire _325_ ;
wire \pp[7]  ;
wire _134_ ;
wire _172_ ;
wire _228_ ;
wire _037_ ;
wire _266_ ;
wire _075_ ;
wire _169_ ;
wire _322_ ;
wire _131_ ;
wire _225_ ;
wire _034_ ;
wire \csa0.y  ;
wire _263_ ;
wire _319_ ;
wire _072_ ;
wire _128_ ;
wire _166_ ;
wire \pp[25]  ;
wire _069_ ;
wire _298_ ;
wire _222_ ;
wire _031_ ;
wire _260_ ;
wire _316_ ;
wire _125_ ;
wire _163_ ;
wire _219_ ;
wire _028_ ;
wire _257_ ;
wire _066_ ;
wire \pp[15]  ;
wire _295_ ;
wire _198_ ;
wire \pp[2]  ;
wire _313_ ;
wire _122_ ;
wire _160_ ;
wire _216_ ;
wire \pp[30]  ;
wire _025_ ;
wire _254_ ;
wire \tcmp.z  ;
wire _063_ ;
wire _119_ ;
wire _292_ ;
wire _157_ ;
wire _195_ ;
wire _289_ ;
wire _098_ ;
wire _310_ ;
wire _213_ ;
wire _022_ ;
wire _251_ ;
wire _307_ ;
wire _060_ ;
wire _116_ ;
wire \pp[20]  ;
wire \pp[9]  ;
wire _154_ ;
wire _019_ ;
wire _192_ ;
wire _248_ ;
wire _057_ ;
wire _286_ ;
wire _095_ ;
wire _189_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _151_ ;
wire _207_ ;
wire _016_ ;
wire \pp[10]  ;
wire _245_ ;
wire _054_ ;
wire _283_ ;
wire _092_ ;
wire _148_ ;
wire _186_ ;
wire \pp[27]  ;
wire _089_ ;
wire _301_ ;
wire _110_ ;
wire _204_ ;
wire _013_ ;
wire _242_ ;
wire _051_ ;
wire _107_ ;
wire _280_ ;
wire _145_ ;
wire _183_ ;
wire _239_ ;
wire _048_ ;
wire _277_ ;
wire _086_ ;
wire \pp[17]  ;
wire _201_ ;
wire _010_ ;
wire \pp[4]  ;
wire _104_ ;
wire _142_ ;
wire _007_ ;
wire _180_ ;
wire _236_ ;
wire _045_ ;
wire _274_ ;
wire _083_ ;
wire _139_ ;
wire _177_ ;
wire _101_ ;
wire _330_ ;
wire _004_ ;
wire _233_ ;
wire _042_ ;
wire _271_ ;
wire _327_ ;
wire _080_ ;
wire _136_ ;
wire \pp[22]  ;
wire _174_ ;
wire _039_ ;
wire _268_ ;
wire _077_ ;
wire clk_1_0 ;
wire _001_ ;
wire _230_ ;
wire _324_ ;
wire _133_ ;
wire _171_ ;
wire _227_ ;
wire _036_ ;
wire \pp[12]  ;
wire _265_ ;
wire _074_ ;

scs8hd_and2_4 _331_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[28]),
    .X(_318_)
);

scs8hd_buf_1 _332_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_318_),
    .X(_319_)
);

scs8hd_o22a_4 _333_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_317_),
    .A1(_316_),
    .X(_320_),
    .B1(_082_),
    .B2(\pp[29] )
);

scs8hd_a2bb2o_4 _334_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_317_),
    .A1N(_316_),
    .X(_038_),
    .B2(_320_),
    .B1(_319_)
);

scs8hd_xor2_4 _335_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_319_),
    .B(_320_),
    .X(_039_)
);

scs8hd_inv_8 _336_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_321_),
    .A(_083_)
);

scs8hd_inv_8 _337_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_322_),
    .A(\pp[30] )
);

scs8hd_and2_4 _338_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[29]),
    .X(_323_)
);

scs8hd_buf_1 _339_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_323_),
    .X(_324_)
);

scs8hd_o22a_4 _340_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_322_),
    .A1(_321_),
    .X(_325_),
    .B1(_083_),
    .B2(\pp[30] )
);

scs8hd_a2bb2o_4 _341_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_322_),
    .A1N(_321_),
    .X(_040_),
    .B2(_325_),
    .B1(_324_)
);

scs8hd_xor2_4 _342_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_324_),
    .B(_325_),
    .X(_041_)
);

scs8hd_inv_8 _343_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_326_),
    .A(_085_)
);

scs8hd_inv_8 _344_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_327_),
    .A(\tcmp.s )
);

scs8hd_and2_4 _345_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .B(x[30]),
    .X(_328_)
);

scs8hd_buf_1 _346_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_328_),
    .X(_329_)
);

scs8hd_o22a_4 _347_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_327_),
    .A1(_326_),
    .X(_330_),
    .B1(_085_),
    .B2(\tcmp.s )
);

scs8hd_a2bb2o_4 _348_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_327_),
    .A1N(_326_),
    .X(_044_),
    .B2(_330_),
    .B1(_329_)
);

scs8hd_xor2_4 _349_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_329_),
    .B(_330_),
    .X(_045_)
);

scs8hd_buf_1 _350_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_156_)
);

scs8hd_inv_8 _351_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_157_),
    .A(rst)
);

scs8hd_buf_1 _352_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_157_),
    .X(_155_)
);

scs8hd_buf_1 _353_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_155_),
    .X(_154_)
);

scs8hd_buf_1 _354_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_155_),
    .X(_153_)
);

scs8hd_buf_1 _355_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_155_),
    .X(_152_)
);

scs8hd_buf_1 _356_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_155_),
    .X(_151_)
);

scs8hd_buf_1 _357_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_155_),
    .X(_150_)
);

scs8hd_buf_1 _358_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_157_),
    .X(_158_)
);

scs8hd_buf_1 _359_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_159_)
);

scs8hd_buf_1 _360_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_149_)
);

scs8hd_buf_1 _361_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_148_)
);

scs8hd_buf_1 _362_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_147_)
);

scs8hd_buf_1 _363_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_146_)
);

scs8hd_buf_1 _364_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_145_)
);

scs8hd_buf_1 _365_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_159_),
    .X(_144_)
);

scs8hd_buf_1 _366_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_160_)
);

scs8hd_buf_1 _367_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_143_)
);

scs8hd_buf_1 _368_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_142_)
);

scs8hd_buf_1 _369_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_141_)
);

scs8hd_buf_1 _370_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_140_)
);

scs8hd_buf_1 _371_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_139_)
);

scs8hd_buf_1 _372_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_160_),
    .X(_138_)
);

scs8hd_buf_1 _373_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_157_),
    .X(_161_)
);

scs8hd_buf_1 _374_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_162_)
);

scs8hd_buf_1 _375_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_137_)
);

scs8hd_buf_1 _376_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_136_)
);

scs8hd_buf_1 _377_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_135_)
);

scs8hd_buf_1 _378_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_134_)
);

scs8hd_buf_1 _379_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_133_)
);

scs8hd_buf_1 _380_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_162_),
    .X(_132_)
);

scs8hd_buf_1 _381_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_163_)
);

scs8hd_buf_1 _382_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_131_)
);

scs8hd_buf_1 _383_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_130_)
);

scs8hd_buf_1 _384_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_129_)
);

scs8hd_buf_1 _385_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_128_)
);

scs8hd_buf_1 _386_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_127_)
);

scs8hd_buf_1 _387_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_163_),
    .X(_126_)
);

scs8hd_buf_1 _388_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_164_)
);

scs8hd_buf_1 _389_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_125_)
);

scs8hd_buf_1 _390_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_124_)
);

scs8hd_buf_1 _391_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_123_)
);

scs8hd_buf_1 _392_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_122_)
);

scs8hd_buf_1 _393_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_121_)
);

scs8hd_buf_1 _394_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_164_),
    .X(_120_)
);

scs8hd_buf_1 _395_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_165_)
);

scs8hd_buf_1 _396_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_119_)
);

scs8hd_buf_1 _397_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_118_)
);

scs8hd_buf_1 _398_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_117_)
);

scs8hd_buf_1 _399_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_116_)
);

scs8hd_buf_1 _400_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_115_)
);

scs8hd_buf_1 _401_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_165_),
    .X(_114_)
);

scs8hd_buf_1 _402_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_166_)
);

scs8hd_buf_1 _403_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_113_)
);

scs8hd_buf_1 _404_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_112_)
);

scs8hd_buf_1 _405_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_111_)
);

scs8hd_buf_1 _406_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_110_)
);

scs8hd_buf_1 _407_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_109_)
);

scs8hd_buf_1 _408_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_166_),
    .X(_108_)
);

scs8hd_buf_1 _409_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_161_),
    .X(_167_)
);

scs8hd_buf_1 _410_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_107_)
);

scs8hd_buf_1 _411_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_106_)
);

scs8hd_buf_1 _412_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_105_)
);

scs8hd_buf_1 _413_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_104_)
);

scs8hd_buf_1 _414_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_103_)
);

scs8hd_buf_1 _415_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_167_),
    .X(_102_)
);

scs8hd_buf_1 _416_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_157_),
    .X(_168_)
);

scs8hd_buf_1 _417_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_101_)
);

scs8hd_buf_1 _418_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_100_)
);

scs8hd_buf_1 _419_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_099_)
);

scs8hd_buf_1 _420_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_098_)
);

scs8hd_buf_1 _421_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_097_)
);

scs8hd_buf_1 _422_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_168_),
    .X(_096_)
);

scs8hd_buf_1 _423_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_095_)
);

scs8hd_buf_1 _424_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_094_)
);

scs8hd_buf_1 _425_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_158_),
    .X(_093_)
);

scs8hd_inv_8 _426_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_169_),
    .A(\csa0.sc )
);

scs8hd_inv_8 _427_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_170_),
    .A(\csa0.y )
);

scs8hd_buf_1 _428_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(y),
    .X(_171_)
);

scs8hd_buf_1 _429_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .X(_172_)
);

scs8hd_and2_4 _430_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[0]),
    .X(_173_)
);

scs8hd_buf_1 _431_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_173_),
    .X(_174_)
);

scs8hd_o22a_4 _432_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_170_),
    .A1(_169_),
    .X(_175_),
    .B1(\csa0.sc ),
    .B2(\csa0.y )
);

scs8hd_a2bb2o_4 _433_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_170_),
    .A1N(_169_),
    .X(_060_),
    .B2(_175_),
    .B1(_174_)
);

scs8hd_xor2_4 _434_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_174_),
    .B(_175_),
    .X(\csa0.hsum2 )
);

scs8hd_and2_4 _435_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .B(x[31]),
    .X(_176_)
);

scs8hd_or2_4 _436_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .B(_176_),
    .A(\tcmp.z ),
    .X(_062_)
);

scs8hd_a21boi_4 _437_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_176_),
    .B1N(_062_),
    .A1(\tcmp.z ),
    .Y(_061_)
);

scs8hd_inv_8 _438_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_177_),
    .A(_073_)
);

scs8hd_inv_8 _439_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_178_),
    .A(\pp[2] )
);

scs8hd_and2_4 _440_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[1]),
    .X(_179_)
);

scs8hd_buf_1 _441_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_179_),
    .X(_180_)
);

scs8hd_o22a_4 _442_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_178_),
    .A1(_177_),
    .X(_181_),
    .B1(_073_),
    .B2(\pp[2] )
);

scs8hd_a2bb2o_4 _443_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_178_),
    .A1N(_177_),
    .X(_020_),
    .B2(_181_),
    .B1(_180_)
);

scs8hd_xor2_4 _444_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_180_),
    .B(_181_),
    .X(_021_)
);

scs8hd_inv_8 _445_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_182_),
    .A(_084_)
);

scs8hd_inv_8 _446_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_183_),
    .A(\pp[3] )
);

scs8hd_and2_4 _447_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[2]),
    .X(_184_)
);

scs8hd_buf_1 _448_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_184_),
    .X(_185_)
);

scs8hd_o22a_4 _449_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_183_),
    .A1(_182_),
    .X(_186_),
    .B1(_084_),
    .B2(\pp[3] )
);

scs8hd_a2bb2o_4 _450_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_183_),
    .A1N(_182_),
    .X(_042_),
    .B2(_186_),
    .B1(_185_)
);

scs8hd_xor2_4 _451_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_185_),
    .B(_186_),
    .X(_043_)
);

scs8hd_inv_8 _452_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_187_),
    .A(_086_)
);

scs8hd_inv_8 _453_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_188_),
    .A(\pp[4] )
);

scs8hd_and2_4 _454_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[3]),
    .X(_189_)
);

scs8hd_buf_1 _455_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_189_),
    .X(_190_)
);

scs8hd_o22a_4 _456_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_188_),
    .A1(_187_),
    .X(_191_),
    .B1(_086_),
    .B2(\pp[4] )
);

scs8hd_a2bb2o_4 _457_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_188_),
    .A1N(_187_),
    .X(_046_),
    .B2(_191_),
    .B1(_190_)
);

scs8hd_xor2_4 _458_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_190_),
    .B(_191_),
    .X(_047_)
);

scs8hd_inv_8 _459_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_192_),
    .A(_087_)
);

scs8hd_inv_8 _460_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_193_),
    .A(\pp[5] )
);

scs8hd_and2_4 _461_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[4]),
    .X(_194_)
);

scs8hd_buf_1 _462_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_194_),
    .X(_195_)
);

scs8hd_o22a_4 _463_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_193_),
    .A1(_192_),
    .X(_196_),
    .B1(_087_),
    .B2(\pp[5] )
);

scs8hd_a2bb2o_4 _464_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_193_),
    .A1N(_192_),
    .X(_048_),
    .B2(_196_),
    .B1(_195_)
);

scs8hd_xor2_4 _465_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_195_),
    .B(_196_),
    .X(_049_)
);

scs8hd_inv_8 _466_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_197_),
    .A(_088_)
);

scs8hd_inv_8 _467_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_198_),
    .A(\pp[6] )
);

scs8hd_and2_4 _468_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_172_),
    .B(x[5]),
    .X(_199_)
);

scs8hd_buf_1 _469_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_199_),
    .X(_200_)
);

scs8hd_o22a_4 _470_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_198_),
    .A1(_197_),
    .X(_201_),
    .B1(_088_),
    .B2(\pp[6] )
);

scs8hd_a2bb2o_4 _471_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_198_),
    .A1N(_197_),
    .X(_050_),
    .B2(_201_),
    .B1(_200_)
);

scs8hd_xor2_4 _472_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_200_),
    .B(_201_),
    .X(_051_)
);

scs8hd_inv_8 _473_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_202_),
    .A(_089_)
);

scs8hd_inv_8 _474_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_203_),
    .A(\pp[7] )
);

scs8hd_buf_1 _475_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .X(_204_)
);

scs8hd_and2_4 _476_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[6]),
    .X(_205_)
);

scs8hd_buf_1 _477_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_205_),
    .X(_206_)
);

scs8hd_o22a_4 _478_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_203_),
    .A1(_202_),
    .X(_207_),
    .B1(_089_),
    .B2(\pp[7] )
);

scs8hd_a2bb2o_4 _479_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_203_),
    .A1N(_202_),
    .X(_052_),
    .B2(_207_),
    .B1(_206_)
);

scs8hd_xor2_4 _480_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_206_),
    .B(_207_),
    .X(_053_)
);

scs8hd_inv_8 _481_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_208_),
    .A(_090_)
);

scs8hd_inv_8 _482_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_209_),
    .A(\pp[8] )
);

scs8hd_and2_4 _483_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[7]),
    .X(_210_)
);

scs8hd_buf_1 _484_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_210_),
    .X(_211_)
);

scs8hd_o22a_4 _485_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_209_),
    .A1(_208_),
    .X(_212_),
    .B1(_090_),
    .B2(\pp[8] )
);

scs8hd_a2bb2o_4 _486_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_209_),
    .A1N(_208_),
    .X(_054_),
    .B2(_212_),
    .B1(_211_)
);

scs8hd_xor2_4 _487_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_211_),
    .B(_212_),
    .X(_055_)
);

scs8hd_inv_8 _488_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_213_),
    .A(_091_)
);

scs8hd_inv_8 _489_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_214_),
    .A(\pp[9] )
);

scs8hd_and2_4 _490_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[8]),
    .X(_215_)
);

scs8hd_buf_1 _491_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_215_),
    .X(_216_)
);

scs8hd_o22a_4 _492_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_214_),
    .A1(_213_),
    .X(_217_),
    .B1(_091_),
    .B2(\pp[9] )
);

scs8hd_a2bb2o_4 _493_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_214_),
    .A1N(_213_),
    .X(_056_),
    .B2(_217_),
    .B1(_216_)
);

scs8hd_xor2_4 _494_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_216_),
    .B(_217_),
    .X(_057_)
);

scs8hd_inv_8 _495_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_218_),
    .A(_092_)
);

scs8hd_inv_8 _496_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_219_),
    .A(\pp[10] )
);

scs8hd_and2_4 _497_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[9]),
    .X(_220_)
);

scs8hd_buf_1 _498_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_220_),
    .X(_221_)
);

scs8hd_o22a_4 _499_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_219_),
    .A1(_218_),
    .X(_222_),
    .B1(_092_),
    .B2(\pp[10] )
);

scs8hd_a2bb2o_4 _500_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_219_),
    .A1N(_218_),
    .X(_058_),
    .B2(_222_),
    .B1(_221_)
);

scs8hd_xor2_4 _501_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_221_),
    .B(_222_),
    .X(_059_)
);

scs8hd_inv_8 _502_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_223_),
    .A(_063_)
);

scs8hd_inv_8 _503_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_224_),
    .A(\pp[11] )
);

scs8hd_and2_4 _504_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[10]),
    .X(_225_)
);

scs8hd_buf_1 _505_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_225_),
    .X(_226_)
);

scs8hd_o22a_4 _506_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_224_),
    .A1(_223_),
    .X(_227_),
    .B1(_063_),
    .B2(\pp[11] )
);

scs8hd_a2bb2o_4 _507_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_224_),
    .A1N(_223_),
    .X(_000_),
    .B2(_227_),
    .B1(_226_)
);

scs8hd_xor2_4 _508_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_226_),
    .B(_227_),
    .X(_001_)
);

scs8hd_inv_8 _509_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_228_),
    .A(_064_)
);

scs8hd_inv_8 _510_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_229_),
    .A(\pp[12] )
);

scs8hd_and2_4 _511_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_204_),
    .B(x[11]),
    .X(_230_)
);

scs8hd_buf_1 _512_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_230_),
    .X(_231_)
);

scs8hd_o22a_4 _513_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_229_),
    .A1(_228_),
    .X(_232_),
    .B1(_064_),
    .B2(\pp[12] )
);

scs8hd_a2bb2o_4 _514_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_229_),
    .A1N(_228_),
    .X(_002_),
    .B2(_232_),
    .B1(_231_)
);

scs8hd_xor2_4 _515_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_231_),
    .B(_232_),
    .X(_003_)
);

scs8hd_inv_8 _516_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_233_),
    .A(_065_)
);

scs8hd_inv_8 _517_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_234_),
    .A(\pp[13] )
);

scs8hd_buf_1 _518_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .X(_235_)
);

scs8hd_and2_4 _519_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[12]),
    .X(_236_)
);

scs8hd_buf_1 _520_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_236_),
    .X(_237_)
);

scs8hd_o22a_4 _521_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_234_),
    .A1(_233_),
    .X(_238_),
    .B1(_065_),
    .B2(\pp[13] )
);

scs8hd_a2bb2o_4 _522_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_234_),
    .A1N(_233_),
    .X(_004_),
    .B2(_238_),
    .B1(_237_)
);

scs8hd_xor2_4 _523_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_237_),
    .B(_238_),
    .X(_005_)
);

scs8hd_inv_8 _524_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_239_),
    .A(_066_)
);

scs8hd_inv_8 _525_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_240_),
    .A(\pp[14] )
);

scs8hd_and2_4 _526_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[13]),
    .X(_241_)
);

scs8hd_buf_1 _527_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_241_),
    .X(_242_)
);

scs8hd_o22a_4 _528_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_240_),
    .A1(_239_),
    .X(_243_),
    .B1(_066_),
    .B2(\pp[14] )
);

scs8hd_a2bb2o_4 _529_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_240_),
    .A1N(_239_),
    .X(_006_),
    .B2(_243_),
    .B1(_242_)
);

scs8hd_xor2_4 _530_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_242_),
    .B(_243_),
    .X(_007_)
);

scs8hd_inv_8 _531_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_244_),
    .A(_067_)
);

scs8hd_inv_8 _532_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_245_),
    .A(\pp[15] )
);

scs8hd_and2_4 _533_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[14]),
    .X(_246_)
);

scs8hd_buf_1 _534_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_246_),
    .X(_247_)
);

scs8hd_o22a_4 _535_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_245_),
    .A1(_244_),
    .X(_248_),
    .B1(_067_),
    .B2(\pp[15] )
);

scs8hd_a2bb2o_4 _536_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_245_),
    .A1N(_244_),
    .X(_008_),
    .B2(_248_),
    .B1(_247_)
);

scs8hd_xor2_4 _537_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_247_),
    .B(_248_),
    .X(_009_)
);

scs8hd_inv_8 _538_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_249_),
    .A(_068_)
);

scs8hd_inv_8 _539_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_250_),
    .A(\pp[16] )
);

scs8hd_and2_4 _540_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[15]),
    .X(_251_)
);

scs8hd_buf_1 _541_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_251_),
    .X(_252_)
);

scs8hd_o22a_4 _542_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_250_),
    .A1(_249_),
    .X(_253_),
    .B1(_068_),
    .B2(\pp[16] )
);

scs8hd_a2bb2o_4 _543_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_250_),
    .A1N(_249_),
    .X(_010_),
    .B2(_253_),
    .B1(_252_)
);

scs8hd_xor2_4 _544_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_252_),
    .B(_253_),
    .X(_011_)
);

scs8hd_inv_8 _545_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_254_),
    .A(_069_)
);

scs8hd_inv_8 _546_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_255_),
    .A(\pp[17] )
);

scs8hd_and2_4 _547_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[16]),
    .X(_256_)
);

scs8hd_buf_1 _548_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_256_),
    .X(_257_)
);

scs8hd_o22a_4 _549_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_255_),
    .A1(_254_),
    .X(_258_),
    .B1(_069_),
    .B2(\pp[17] )
);

scs8hd_a2bb2o_4 _550_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_255_),
    .A1N(_254_),
    .X(_012_),
    .B2(_258_),
    .B1(_257_)
);

scs8hd_xor2_4 _551_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_257_),
    .B(_258_),
    .X(_013_)
);

scs8hd_inv_8 _552_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_259_),
    .A(_070_)
);

scs8hd_inv_8 _553_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_260_),
    .A(\pp[18] )
);

scs8hd_and2_4 _554_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_235_),
    .B(x[17]),
    .X(_261_)
);

scs8hd_buf_1 _555_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_261_),
    .X(_262_)
);

scs8hd_o22a_4 _556_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_260_),
    .A1(_259_),
    .X(_263_),
    .B1(_070_),
    .B2(\pp[18] )
);

scs8hd_a2bb2o_4 _557_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_260_),
    .A1N(_259_),
    .X(_014_),
    .B2(_263_),
    .B1(_262_)
);

scs8hd_xor2_4 _558_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_262_),
    .B(_263_),
    .X(_015_)
);

scs8hd_inv_8 _559_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_264_),
    .A(_071_)
);

scs8hd_inv_8 _560_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_265_),
    .A(\pp[19] )
);

scs8hd_buf_1 _561_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_171_),
    .X(_266_)
);

scs8hd_and2_4 _562_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[18]),
    .X(_267_)
);

scs8hd_buf_1 _563_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_267_),
    .X(_268_)
);

scs8hd_o22a_4 _564_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_265_),
    .A1(_264_),
    .X(_269_),
    .B1(_071_),
    .B2(\pp[19] )
);

scs8hd_a2bb2o_4 _565_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_265_),
    .A1N(_264_),
    .X(_016_),
    .B2(_269_),
    .B1(_268_)
);

scs8hd_xor2_4 _566_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_268_),
    .B(_269_),
    .X(_017_)
);

scs8hd_inv_8 _567_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_270_),
    .A(_072_)
);

scs8hd_inv_8 _568_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_271_),
    .A(\pp[20] )
);

scs8hd_and2_4 _569_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[19]),
    .X(_272_)
);

scs8hd_buf_1 _570_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_272_),
    .X(_273_)
);

scs8hd_o22a_4 _571_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_271_),
    .A1(_270_),
    .X(_274_),
    .B1(_072_),
    .B2(\pp[20] )
);

scs8hd_a2bb2o_4 _572_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_271_),
    .A1N(_270_),
    .X(_018_),
    .B2(_274_),
    .B1(_273_)
);

scs8hd_xor2_4 _573_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_273_),
    .B(_274_),
    .X(_019_)
);

scs8hd_inv_8 _574_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_275_),
    .A(_074_)
);

scs8hd_inv_8 _575_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_276_),
    .A(\pp[21] )
);

scs8hd_and2_4 _576_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[20]),
    .X(_277_)
);

scs8hd_buf_1 _577_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_277_),
    .X(_278_)
);

scs8hd_o22a_4 _578_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_276_),
    .A1(_275_),
    .X(_279_),
    .B1(_074_),
    .B2(\pp[21] )
);

scs8hd_a2bb2o_4 _579_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_276_),
    .A1N(_275_),
    .X(_022_),
    .B2(_279_),
    .B1(_278_)
);

scs8hd_xor2_4 _580_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_278_),
    .B(_279_),
    .X(_023_)
);

scs8hd_inv_8 _581_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_280_),
    .A(_075_)
);

scs8hd_inv_8 _582_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_281_),
    .A(\pp[22] )
);

scs8hd_and2_4 _583_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[21]),
    .X(_282_)
);

scs8hd_buf_1 _584_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_282_),
    .X(_283_)
);

scs8hd_o22a_4 _585_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_281_),
    .A1(_280_),
    .X(_284_),
    .B1(_075_),
    .B2(\pp[22] )
);

scs8hd_a2bb2o_4 _586_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_281_),
    .A1N(_280_),
    .X(_024_),
    .B2(_284_),
    .B1(_283_)
);

scs8hd_xor2_4 _587_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_283_),
    .B(_284_),
    .X(_025_)
);

scs8hd_inv_8 _588_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_285_),
    .A(_076_)
);

scs8hd_inv_8 _589_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_286_),
    .A(\pp[23] )
);

scs8hd_and2_4 _590_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[22]),
    .X(_287_)
);

scs8hd_buf_1 _591_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_287_),
    .X(_288_)
);

scs8hd_o22a_4 _592_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_286_),
    .A1(_285_),
    .X(_289_),
    .B1(_076_),
    .B2(\pp[23] )
);

scs8hd_a2bb2o_4 _593_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_286_),
    .A1N(_285_),
    .X(_026_),
    .B2(_289_),
    .B1(_288_)
);

scs8hd_xor2_4 _594_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_288_),
    .B(_289_),
    .X(_027_)
);

scs8hd_inv_8 _595_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_290_),
    .A(_077_)
);

scs8hd_inv_8 _596_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_291_),
    .A(\pp[24] )
);

scs8hd_and2_4 _597_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_266_),
    .B(x[23]),
    .X(_292_)
);

scs8hd_buf_1 _598_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_292_),
    .X(_293_)
);

scs8hd_o22a_4 _599_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_291_),
    .A1(_290_),
    .X(_294_),
    .B1(_077_),
    .B2(\pp[24] )
);

scs8hd_a2bb2o_4 _600_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_291_),
    .A1N(_290_),
    .X(_028_),
    .B2(_294_),
    .B1(_293_)
);

scs8hd_xor2_4 _601_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_293_),
    .B(_294_),
    .X(_029_)
);

scs8hd_inv_8 _602_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_295_),
    .A(_078_)
);

scs8hd_inv_8 _603_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_296_),
    .A(\pp[25] )
);

scs8hd_buf_1 _604_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(y),
    .X(_297_)
);

scs8hd_and2_4 _605_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[24]),
    .X(_298_)
);

scs8hd_buf_1 _606_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_298_),
    .X(_299_)
);

scs8hd_o22a_4 _607_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_296_),
    .A1(_295_),
    .X(_300_),
    .B1(_078_),
    .B2(\pp[25] )
);

scs8hd_a2bb2o_4 _608_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_296_),
    .A1N(_295_),
    .X(_030_),
    .B2(_300_),
    .B1(_299_)
);

scs8hd_xor2_4 _609_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_299_),
    .B(_300_),
    .X(_031_)
);

scs8hd_inv_8 _610_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_301_),
    .A(_079_)
);

scs8hd_inv_8 _611_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_302_),
    .A(\pp[26] )
);

scs8hd_and2_4 _612_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[25]),
    .X(_303_)
);

scs8hd_buf_1 _613_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_303_),
    .X(_304_)
);

scs8hd_o22a_4 _614_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_302_),
    .A1(_301_),
    .X(_305_),
    .B1(_079_),
    .B2(\pp[26] )
);

scs8hd_a2bb2o_4 _615_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_302_),
    .A1N(_301_),
    .X(_032_),
    .B2(_305_),
    .B1(_304_)
);

scs8hd_xor2_4 _616_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_304_),
    .B(_305_),
    .X(_033_)
);

scs8hd_inv_8 _617_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_306_),
    .A(_080_)
);

scs8hd_inv_8 _618_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_307_),
    .A(\pp[27] )
);

scs8hd_and2_4 _619_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[26]),
    .X(_308_)
);

scs8hd_buf_1 _620_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_308_),
    .X(_309_)
);

scs8hd_o22a_4 _621_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_307_),
    .A1(_306_),
    .X(_310_),
    .B1(_080_),
    .B2(\pp[27] )
);

scs8hd_a2bb2o_4 _622_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_307_),
    .A1N(_306_),
    .X(_034_),
    .B2(_310_),
    .B1(_309_)
);

scs8hd_xor2_4 _623_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_309_),
    .B(_310_),
    .X(_035_)
);

scs8hd_inv_8 _624_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_311_),
    .A(_081_)
);

scs8hd_inv_8 _625_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_312_),
    .A(\pp[28] )
);

scs8hd_and2_4 _626_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_297_),
    .B(x[27]),
    .X(_313_)
);

scs8hd_buf_1 _627_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_313_),
    .X(_314_)
);

scs8hd_o22a_4 _628_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2(_312_),
    .A1(_311_),
    .X(_315_),
    .B1(_081_),
    .B2(\pp[28] )
);

scs8hd_a2bb2o_4 _629_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A2N(_312_),
    .A1N(_311_),
    .X(_036_),
    .B2(_315_),
    .B1(_314_)
);

scs8hd_xor2_4 _630_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(_314_),
    .B(_315_),
    .X(_037_)
);

scs8hd_inv_8 _631_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_316_),
    .A(_082_)
);

scs8hd_inv_8 _632_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .Y(_317_),
    .A(\pp[29] )
);

scs8hd_dfrtp_4 _633_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_060_),
    .RESETB(_093_),
    .Q(\csa0.sc )
);

scs8hd_dfrtp_4 _634_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(\csa0.hsum2 ),
    .RESETB(_094_),
    .Q(p)
);

scs8hd_dfrtp_4 _635_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_062_),
    .RESETB(_095_),
    .Q(\tcmp.z )
);

scs8hd_dfrtp_4 _636_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_061_),
    .RESETB(_096_),
    .Q(\tcmp.s )
);

scs8hd_dfrtp_4 _637_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_020_),
    .RESETB(_097_),
    .Q(_073_)
);

scs8hd_dfrtp_4 _638_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_021_),
    .RESETB(_098_),
    .Q(\csa0.y )
);

scs8hd_dfrtp_4 _639_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_042_),
    .RESETB(_099_),
    .Q(_084_)
);

scs8hd_dfrtp_4 _640_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_043_),
    .RESETB(_100_),
    .Q(\pp[2] )
);

scs8hd_dfrtp_4 _641_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_046_),
    .RESETB(_101_),
    .Q(_086_)
);

scs8hd_dfrtp_4 _642_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_047_),
    .RESETB(_102_),
    .Q(\pp[3] )
);

scs8hd_dfrtp_4 _643_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_048_),
    .RESETB(_103_),
    .Q(_087_)
);

scs8hd_dfrtp_4 _644_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_049_),
    .RESETB(_104_),
    .Q(\pp[4] )
);

scs8hd_dfrtp_4 _645_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_050_),
    .RESETB(_105_),
    .Q(_088_)
);

scs8hd_dfrtp_4 _646_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_051_),
    .RESETB(_106_),
    .Q(\pp[5] )
);

scs8hd_dfrtp_4 _647_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_052_),
    .RESETB(_107_),
    .Q(_089_)
);

scs8hd_dfrtp_4 _648_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_0),
    .D(_053_),
    .RESETB(_108_),
    .Q(\pp[6] )
);

scs8hd_dfrtp_4 _649_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_054_),
    .RESETB(_109_),
    .Q(_090_)
);

scs8hd_dfrtp_4 _650_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_055_),
    .RESETB(_110_),
    .Q(\pp[7] )
);

scs8hd_dfrtp_4 _651_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_056_),
    .RESETB(_111_),
    .Q(_091_)
);

scs8hd_dfrtp_4 _652_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_057_),
    .RESETB(_112_),
    .Q(\pp[8] )
);

scs8hd_dfrtp_4 _653_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_058_),
    .RESETB(_113_),
    .Q(_092_)
);

scs8hd_dfrtp_4 _654_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_059_),
    .RESETB(_114_),
    .Q(\pp[9] )
);

scs8hd_dfrtp_4 _655_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_000_),
    .RESETB(_115_),
    .Q(_063_)
);

scs8hd_dfrtp_4 _656_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_001_),
    .RESETB(_116_),
    .Q(\pp[10] )
);

scs8hd_dfrtp_4 _657_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_002_),
    .RESETB(_117_),
    .Q(_064_)
);

scs8hd_dfrtp_4 _658_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_003_),
    .RESETB(_118_),
    .Q(\pp[11] )
);

scs8hd_dfrtp_4 _659_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_004_),
    .RESETB(_119_),
    .Q(_065_)
);

scs8hd_dfrtp_4 _660_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_005_),
    .RESETB(_120_),
    .Q(\pp[12] )
);

scs8hd_dfrtp_4 _661_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_006_),
    .RESETB(_121_),
    .Q(_066_)
);

scs8hd_dfrtp_4 _662_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_007_),
    .RESETB(_122_),
    .Q(\pp[13] )
);

scs8hd_dfrtp_4 _663_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_008_),
    .RESETB(_123_),
    .Q(_067_)
);

scs8hd_dfrtp_4 _664_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_16),
    .D(_009_),
    .RESETB(_124_),
    .Q(\pp[14] )
);

scs8hd_dfrtp_4 _665_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_010_),
    .RESETB(_125_),
    .Q(_068_)
);

scs8hd_dfrtp_4 _666_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_011_),
    .RESETB(_126_),
    .Q(\pp[15] )
);

scs8hd_dfrtp_4 _667_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_012_),
    .RESETB(_127_),
    .Q(_069_)
);

scs8hd_dfrtp_4 _668_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_013_),
    .RESETB(_128_),
    .Q(\pp[16] )
);

scs8hd_dfrtp_4 _669_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_014_),
    .RESETB(_129_),
    .Q(_070_)
);

scs8hd_dfrtp_4 _670_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_015_),
    .RESETB(_130_),
    .Q(\pp[17] )
);

scs8hd_dfrtp_4 _671_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_016_),
    .RESETB(_131_),
    .Q(_071_)
);

scs8hd_dfrtp_4 _672_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_017_),
    .RESETB(_132_),
    .Q(\pp[18] )
);

scs8hd_dfrtp_4 _673_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_018_),
    .RESETB(_133_),
    .Q(_072_)
);

scs8hd_dfrtp_4 _674_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_019_),
    .RESETB(_134_),
    .Q(\pp[19] )
);

scs8hd_dfrtp_4 _675_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_022_),
    .RESETB(_135_),
    .Q(_074_)
);

scs8hd_dfrtp_4 _676_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_023_),
    .RESETB(_136_),
    .Q(\pp[20] )
);

scs8hd_dfrtp_4 _677_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_024_),
    .RESETB(_137_),
    .Q(_075_)
);

scs8hd_dfrtp_4 _678_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_025_),
    .RESETB(_138_),
    .Q(\pp[21] )
);

scs8hd_dfrtp_4 _679_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_026_),
    .RESETB(_139_),
    .Q(_076_)
);

scs8hd_dfrtp_4 _680_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_32),
    .D(_027_),
    .RESETB(_140_),
    .Q(\pp[22] )
);

scs8hd_dfrtp_4 _681_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_028_),
    .RESETB(_141_),
    .Q(_077_)
);

scs8hd_dfrtp_4 _682_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_029_),
    .RESETB(_142_),
    .Q(\pp[23] )
);

scs8hd_dfrtp_4 _683_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_030_),
    .RESETB(_143_),
    .Q(_078_)
);

scs8hd_dfrtp_4 _684_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_031_),
    .RESETB(_144_),
    .Q(\pp[24] )
);

scs8hd_dfrtp_4 _685_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_032_),
    .RESETB(_145_),
    .Q(_079_)
);

scs8hd_dfrtp_4 _686_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_033_),
    .RESETB(_146_),
    .Q(\pp[25] )
);

scs8hd_dfrtp_4 _687_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_034_),
    .RESETB(_147_),
    .Q(_080_)
);

scs8hd_dfrtp_4 _688_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_035_),
    .RESETB(_148_),
    .Q(\pp[26] )
);

scs8hd_dfrtp_4 _689_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_036_),
    .RESETB(_149_),
    .Q(_081_)
);

scs8hd_dfrtp_4 _690_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_037_),
    .RESETB(_150_),
    .Q(\pp[27] )
);

scs8hd_dfrtp_4 _691_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_038_),
    .RESETB(_151_),
    .Q(_082_)
);

scs8hd_dfrtp_4 _692_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_039_),
    .RESETB(_152_),
    .Q(\pp[28] )
);

scs8hd_dfrtp_4 _693_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_040_),
    .RESETB(_153_),
    .Q(_083_)
);

scs8hd_dfrtp_4 _694_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_041_),
    .RESETB(_154_),
    .Q(\pp[29] )
);

scs8hd_dfrtp_4 _695_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_044_),
    .RESETB(_155_),
    .Q(_085_)
);

scs8hd_dfrtp_4 _696_ (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .CLK(clk_0_48),
    .D(_045_),
    .RESETB(_156_),
    .Q(\pp[30] )
);

scs8hd_clkbuf_4 _CTS_buf_1_0 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(clk_1_0),
    .X(clk_0_0)
);

scs8hd_clkbuf_4 _CTS_buf_1_16 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(clk_1_0),
    .X(clk_0_16)
);

scs8hd_clkbuf_4 _CTS_buf_1_32 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(clk_1_0),
    .X(clk_0_32)
);

scs8hd_clkbuf_4 _CTS_buf_1_48 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(clk_1_0),
    .X(clk_0_48)
);

scs8hd_clkbuf_16 _CTS_root (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .A(clk),
    .X(clk_1_0)
);

scs8hd_decap_3 PHY_0 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_1 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_2 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_3 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_4 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_5 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_6 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_7 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_8 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_9 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_10 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_11 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_12 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_13 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_14 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_15 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_16 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_17 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_18 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_19 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_20 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_21 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_22 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_23 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_24 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_25 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_26 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_27 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_28 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_29 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_30 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_31 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_32 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_33 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_34 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_35 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_36 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_37 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_38 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_39 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_40 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_41 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_42 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_43 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_44 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_45 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_46 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_47 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_48 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_49 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_50 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_51 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_52 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_53 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_54 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_55 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_56 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_57 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_58 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_59 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_60 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_61 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_62 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_63 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_64 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_65 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_66 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_67 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_68 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_69 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_70 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_71 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_72 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_73 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_74 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_75 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_76 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_77 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_78 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_79 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_80 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_81 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_82 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_83 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_84 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_decap_3 PHY_85 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_86 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_87 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_88 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_89 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_90 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_91 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_92 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_93 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_94 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_95 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_96 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_97 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_98 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_99 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_100 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_101 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_102 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_103 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_104 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_105 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_106 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_107 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_108 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_109 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_110 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_111 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_112 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_113 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_114 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_115 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_116 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_117 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_118 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_119 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_120 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_121 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_122 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_123 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_124 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_125 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_126 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_127 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_128 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_129 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_130 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_131 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_132 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_133 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_134 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_135 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_136 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_137 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_138 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_139 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_140 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_141 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_142 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_143 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_144 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_145 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_146 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_147 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_148 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_149 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_150 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_151 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_152 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_153 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_154 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_155 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_156 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_157 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_158 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_159 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_160 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_161 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_162 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_163 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_164 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_165 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_166 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_167 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_168 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_169 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_170 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_171 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_172 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_173 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_174 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_175 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_176 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_177 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_178 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_179 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_180 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_181 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_182 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_183 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_184 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_185 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_186 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_187 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_188 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_189 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_190 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_191 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_192 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_193 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_194 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_195 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_196 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_197 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_198 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_199 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_200 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_201 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_202 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_203 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_204 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_205 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_206 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_207 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_208 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_209 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_210 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_211 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_212 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_213 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_214 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_215 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_216 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_217 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_218 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_219 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_220 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_221 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_222 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_223 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_224 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_225 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_226 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_227 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_228 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_229 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_230 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_231 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_232 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_233 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_234 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_235 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_236 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_237 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_238 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_239 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_240 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_241 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_242 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_243 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_244 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_245 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_246 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_247 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_248 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_249 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_250 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_251 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_252 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_253 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_254 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_255 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_256 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_257 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_258 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_259 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_260 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_261 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_262 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_263 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_264 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_tapvpwrvgnd_1 PHY_265 (
    .vgnd(vgnd),
    .vpwr(vpwr)
);

scs8hd_diode_2 ANTENNA__CTS_root_A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk)
);

scs8hd_diode_2 ANTENNA__351__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(rst)
);

scs8hd_diode_2 ANTENNA__430__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[0])
);

scs8hd_diode_2 ANTENNA__504__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[10])
);

scs8hd_diode_2 ANTENNA__511__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[11])
);

scs8hd_diode_2 ANTENNA__519__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[12])
);

scs8hd_diode_2 ANTENNA__526__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[13])
);

scs8hd_diode_2 ANTENNA__533__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[14])
);

scs8hd_diode_2 ANTENNA__540__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[15])
);

scs8hd_diode_2 ANTENNA__547__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[16])
);

scs8hd_diode_2 ANTENNA__554__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[17])
);

scs8hd_diode_2 ANTENNA__562__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[18])
);

scs8hd_diode_2 ANTENNA__569__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[19])
);

scs8hd_diode_2 ANTENNA__440__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[1])
);

scs8hd_diode_2 ANTENNA__576__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[20])
);

scs8hd_diode_2 ANTENNA__583__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[21])
);

scs8hd_diode_2 ANTENNA__590__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[22])
);

scs8hd_diode_2 ANTENNA__597__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[23])
);

scs8hd_diode_2 ANTENNA__605__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[24])
);

scs8hd_diode_2 ANTENNA__612__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[25])
);

scs8hd_diode_2 ANTENNA__619__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[26])
);

scs8hd_diode_2 ANTENNA__626__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[27])
);

scs8hd_diode_2 ANTENNA__331__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[28])
);

scs8hd_diode_2 ANTENNA__338__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[29])
);

scs8hd_diode_2 ANTENNA__447__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[2])
);

scs8hd_diode_2 ANTENNA__345__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[30])
);

scs8hd_diode_2 ANTENNA__435__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[31])
);

scs8hd_diode_2 ANTENNA__454__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[3])
);

scs8hd_diode_2 ANTENNA__461__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[4])
);

scs8hd_diode_2 ANTENNA__468__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[5])
);

scs8hd_diode_2 ANTENNA__476__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[6])
);

scs8hd_diode_2 ANTENNA__483__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[7])
);

scs8hd_diode_2 ANTENNA__490__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[8])
);

scs8hd_diode_2 ANTENNA__497__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(x[9])
);

scs8hd_diode_2 ANTENNA__604__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(y)
);

scs8hd_diode_2 ANTENNA__428__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(y)
);

scs8hd_diode_2 ANTENNA__655__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_000_)
);

scs8hd_diode_2 ANTENNA__656__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_001_)
);

scs8hd_diode_2 ANTENNA__657__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_002_)
);

scs8hd_diode_2 ANTENNA__658__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_003_)
);

scs8hd_diode_2 ANTENNA__659__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_004_)
);

scs8hd_diode_2 ANTENNA__660__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_005_)
);

scs8hd_diode_2 ANTENNA__661__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_006_)
);

scs8hd_diode_2 ANTENNA__662__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_007_)
);

scs8hd_diode_2 ANTENNA__663__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_008_)
);

scs8hd_diode_2 ANTENNA__664__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_009_)
);

scs8hd_diode_2 ANTENNA__665__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_010_)
);

scs8hd_diode_2 ANTENNA__666__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_011_)
);

scs8hd_diode_2 ANTENNA__667__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_012_)
);

scs8hd_diode_2 ANTENNA__668__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_013_)
);

scs8hd_diode_2 ANTENNA__669__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_014_)
);

scs8hd_diode_2 ANTENNA__670__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_015_)
);

scs8hd_diode_2 ANTENNA__671__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_016_)
);

scs8hd_diode_2 ANTENNA__672__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_017_)
);

scs8hd_diode_2 ANTENNA__673__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_018_)
);

scs8hd_diode_2 ANTENNA__674__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_019_)
);

scs8hd_diode_2 ANTENNA__637__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_020_)
);

scs8hd_diode_2 ANTENNA__638__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_021_)
);

scs8hd_diode_2 ANTENNA__675__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_022_)
);

scs8hd_diode_2 ANTENNA__676__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_023_)
);

scs8hd_diode_2 ANTENNA__677__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_024_)
);

scs8hd_diode_2 ANTENNA__678__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_025_)
);

scs8hd_diode_2 ANTENNA__679__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_026_)
);

scs8hd_diode_2 ANTENNA__680__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_027_)
);

scs8hd_diode_2 ANTENNA__681__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_028_)
);

scs8hd_diode_2 ANTENNA__682__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_029_)
);

scs8hd_diode_2 ANTENNA__683__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_030_)
);

scs8hd_diode_2 ANTENNA__684__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_031_)
);

scs8hd_diode_2 ANTENNA__685__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_032_)
);

scs8hd_diode_2 ANTENNA__686__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_033_)
);

scs8hd_diode_2 ANTENNA__687__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_034_)
);

scs8hd_diode_2 ANTENNA__688__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_035_)
);

scs8hd_diode_2 ANTENNA__689__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_036_)
);

scs8hd_diode_2 ANTENNA__690__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_037_)
);

scs8hd_diode_2 ANTENNA__691__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_038_)
);

scs8hd_diode_2 ANTENNA__692__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_039_)
);

scs8hd_diode_2 ANTENNA__693__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_040_)
);

scs8hd_diode_2 ANTENNA__694__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_041_)
);

scs8hd_diode_2 ANTENNA__639__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_042_)
);

scs8hd_diode_2 ANTENNA__640__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_043_)
);

scs8hd_diode_2 ANTENNA__695__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_044_)
);

scs8hd_diode_2 ANTENNA__696__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_045_)
);

scs8hd_diode_2 ANTENNA__641__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_046_)
);

scs8hd_diode_2 ANTENNA__642__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_047_)
);

scs8hd_diode_2 ANTENNA__643__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_048_)
);

scs8hd_diode_2 ANTENNA__644__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_049_)
);

scs8hd_diode_2 ANTENNA__645__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_050_)
);

scs8hd_diode_2 ANTENNA__646__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_051_)
);

scs8hd_diode_2 ANTENNA__647__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_052_)
);

scs8hd_diode_2 ANTENNA__648__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_053_)
);

scs8hd_diode_2 ANTENNA__649__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_054_)
);

scs8hd_diode_2 ANTENNA__650__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_055_)
);

scs8hd_diode_2 ANTENNA__651__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_056_)
);

scs8hd_diode_2 ANTENNA__652__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_057_)
);

scs8hd_diode_2 ANTENNA__653__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_058_)
);

scs8hd_diode_2 ANTENNA__654__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_059_)
);

scs8hd_diode_2 ANTENNA__633__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_060_)
);

scs8hd_diode_2 ANTENNA__636__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_061_)
);

scs8hd_diode_2 ANTENNA__635__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_062_)
);

scs8hd_diode_2 ANTENNA__437__B1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_062_)
);

scs8hd_diode_2 ANTENNA__506__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_063_)
);

scs8hd_diode_2 ANTENNA__502__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_063_)
);

scs8hd_diode_2 ANTENNA__513__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_064_)
);

scs8hd_diode_2 ANTENNA__509__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_064_)
);

scs8hd_diode_2 ANTENNA__521__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_065_)
);

scs8hd_diode_2 ANTENNA__516__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_065_)
);

scs8hd_diode_2 ANTENNA__528__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_066_)
);

scs8hd_diode_2 ANTENNA__524__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_066_)
);

scs8hd_diode_2 ANTENNA__535__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_067_)
);

scs8hd_diode_2 ANTENNA__531__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_067_)
);

scs8hd_diode_2 ANTENNA__542__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_068_)
);

scs8hd_diode_2 ANTENNA__538__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_068_)
);

scs8hd_diode_2 ANTENNA__549__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_069_)
);

scs8hd_diode_2 ANTENNA__545__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_069_)
);

scs8hd_diode_2 ANTENNA__556__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_070_)
);

scs8hd_diode_2 ANTENNA__552__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_070_)
);

scs8hd_diode_2 ANTENNA__564__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_071_)
);

scs8hd_diode_2 ANTENNA__559__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_071_)
);

scs8hd_diode_2 ANTENNA__571__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_072_)
);

scs8hd_diode_2 ANTENNA__567__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_072_)
);

scs8hd_diode_2 ANTENNA__442__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_073_)
);

scs8hd_diode_2 ANTENNA__438__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_073_)
);

scs8hd_diode_2 ANTENNA__578__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_074_)
);

scs8hd_diode_2 ANTENNA__574__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_074_)
);

scs8hd_diode_2 ANTENNA__585__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_075_)
);

scs8hd_diode_2 ANTENNA__581__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_075_)
);

scs8hd_diode_2 ANTENNA__592__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_076_)
);

scs8hd_diode_2 ANTENNA__588__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_076_)
);

scs8hd_diode_2 ANTENNA__599__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_077_)
);

scs8hd_diode_2 ANTENNA__595__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_077_)
);

scs8hd_diode_2 ANTENNA__607__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_078_)
);

scs8hd_diode_2 ANTENNA__602__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_078_)
);

scs8hd_diode_2 ANTENNA__614__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_079_)
);

scs8hd_diode_2 ANTENNA__610__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_079_)
);

scs8hd_diode_2 ANTENNA__621__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_080_)
);

scs8hd_diode_2 ANTENNA__617__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_080_)
);

scs8hd_diode_2 ANTENNA__628__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_081_)
);

scs8hd_diode_2 ANTENNA__624__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_081_)
);

scs8hd_diode_2 ANTENNA__631__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_082_)
);

scs8hd_diode_2 ANTENNA__333__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_082_)
);

scs8hd_diode_2 ANTENNA__340__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_083_)
);

scs8hd_diode_2 ANTENNA__336__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_083_)
);

scs8hd_diode_2 ANTENNA__449__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_084_)
);

scs8hd_diode_2 ANTENNA__445__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_084_)
);

scs8hd_diode_2 ANTENNA__347__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_085_)
);

scs8hd_diode_2 ANTENNA__343__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_085_)
);

scs8hd_diode_2 ANTENNA__456__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_086_)
);

scs8hd_diode_2 ANTENNA__452__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_086_)
);

scs8hd_diode_2 ANTENNA__463__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_087_)
);

scs8hd_diode_2 ANTENNA__459__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_087_)
);

scs8hd_diode_2 ANTENNA__470__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_088_)
);

scs8hd_diode_2 ANTENNA__466__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_088_)
);

scs8hd_diode_2 ANTENNA__478__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_089_)
);

scs8hd_diode_2 ANTENNA__473__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_089_)
);

scs8hd_diode_2 ANTENNA__485__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_090_)
);

scs8hd_diode_2 ANTENNA__481__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_090_)
);

scs8hd_diode_2 ANTENNA__492__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_091_)
);

scs8hd_diode_2 ANTENNA__488__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_091_)
);

scs8hd_diode_2 ANTENNA__499__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_092_)
);

scs8hd_diode_2 ANTENNA__495__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_092_)
);

scs8hd_diode_2 ANTENNA__633__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_093_)
);

scs8hd_diode_2 ANTENNA__634__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_094_)
);

scs8hd_diode_2 ANTENNA__635__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_095_)
);

scs8hd_diode_2 ANTENNA__636__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_096_)
);

scs8hd_diode_2 ANTENNA__637__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_097_)
);

scs8hd_diode_2 ANTENNA__638__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_098_)
);

scs8hd_diode_2 ANTENNA__639__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_099_)
);

scs8hd_diode_2 ANTENNA__640__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_100_)
);

scs8hd_diode_2 ANTENNA__641__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_101_)
);

scs8hd_diode_2 ANTENNA__642__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_102_)
);

scs8hd_diode_2 ANTENNA__643__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_103_)
);

scs8hd_diode_2 ANTENNA__644__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_104_)
);

scs8hd_diode_2 ANTENNA__645__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_105_)
);

scs8hd_diode_2 ANTENNA__646__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_106_)
);

scs8hd_diode_2 ANTENNA__647__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_107_)
);

scs8hd_diode_2 ANTENNA__648__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_108_)
);

scs8hd_diode_2 ANTENNA__649__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_109_)
);

scs8hd_diode_2 ANTENNA__650__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_110_)
);

scs8hd_diode_2 ANTENNA__651__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_111_)
);

scs8hd_diode_2 ANTENNA__652__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_112_)
);

scs8hd_diode_2 ANTENNA__653__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_113_)
);

scs8hd_diode_2 ANTENNA__654__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_114_)
);

scs8hd_diode_2 ANTENNA__655__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_115_)
);

scs8hd_diode_2 ANTENNA__656__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_116_)
);

scs8hd_diode_2 ANTENNA__657__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_117_)
);

scs8hd_diode_2 ANTENNA__658__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_118_)
);

scs8hd_diode_2 ANTENNA__659__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_119_)
);

scs8hd_diode_2 ANTENNA__660__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_120_)
);

scs8hd_diode_2 ANTENNA__661__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_121_)
);

scs8hd_diode_2 ANTENNA__662__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_122_)
);

scs8hd_diode_2 ANTENNA__663__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_123_)
);

scs8hd_diode_2 ANTENNA__664__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_124_)
);

scs8hd_diode_2 ANTENNA__665__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_125_)
);

scs8hd_diode_2 ANTENNA__666__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_126_)
);

scs8hd_diode_2 ANTENNA__667__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_127_)
);

scs8hd_diode_2 ANTENNA__668__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_128_)
);

scs8hd_diode_2 ANTENNA__669__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_129_)
);

scs8hd_diode_2 ANTENNA__670__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_130_)
);

scs8hd_diode_2 ANTENNA__671__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_131_)
);

scs8hd_diode_2 ANTENNA__672__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_132_)
);

scs8hd_diode_2 ANTENNA__673__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_133_)
);

scs8hd_diode_2 ANTENNA__674__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_134_)
);

scs8hd_diode_2 ANTENNA__675__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_135_)
);

scs8hd_diode_2 ANTENNA__676__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_136_)
);

scs8hd_diode_2 ANTENNA__677__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_137_)
);

scs8hd_diode_2 ANTENNA__678__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_138_)
);

scs8hd_diode_2 ANTENNA__679__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_139_)
);

scs8hd_diode_2 ANTENNA__680__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_140_)
);

scs8hd_diode_2 ANTENNA__681__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_141_)
);

scs8hd_diode_2 ANTENNA__682__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_142_)
);

scs8hd_diode_2 ANTENNA__683__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_143_)
);

scs8hd_diode_2 ANTENNA__684__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_144_)
);

scs8hd_diode_2 ANTENNA__685__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_145_)
);

scs8hd_diode_2 ANTENNA__686__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_146_)
);

scs8hd_diode_2 ANTENNA__687__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_147_)
);

scs8hd_diode_2 ANTENNA__688__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_148_)
);

scs8hd_diode_2 ANTENNA__689__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_149_)
);

scs8hd_diode_2 ANTENNA__690__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_150_)
);

scs8hd_diode_2 ANTENNA__691__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_151_)
);

scs8hd_diode_2 ANTENNA__692__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_152_)
);

scs8hd_diode_2 ANTENNA__693__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_153_)
);

scs8hd_diode_2 ANTENNA__694__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_154_)
);

scs8hd_diode_2 ANTENNA__695__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__357__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__356__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__355__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__354__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__353__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_155_)
);

scs8hd_diode_2 ANTENNA__696__RESETB (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_156_)
);

scs8hd_diode_2 ANTENNA__416__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_157_)
);

scs8hd_diode_2 ANTENNA__373__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_157_)
);

scs8hd_diode_2 ANTENNA__358__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_157_)
);

scs8hd_diode_2 ANTENNA__352__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_157_)
);

scs8hd_diode_2 ANTENNA__425__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__424__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__423__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__366__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__359__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__350__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_158_)
);

scs8hd_diode_2 ANTENNA__365__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__364__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__363__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__362__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__361__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__360__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_159_)
);

scs8hd_diode_2 ANTENNA__372__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__371__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__370__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__369__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__368__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__367__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_160_)
);

scs8hd_diode_2 ANTENNA__409__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__402__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__395__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__388__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__381__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__374__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_161_)
);

scs8hd_diode_2 ANTENNA__380__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__379__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__378__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__377__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__376__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__375__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_162_)
);

scs8hd_diode_2 ANTENNA__387__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__386__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__385__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__384__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__383__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__382__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_163_)
);

scs8hd_diode_2 ANTENNA__394__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__393__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__392__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__391__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__390__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__389__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_164_)
);

scs8hd_diode_2 ANTENNA__401__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__400__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__399__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__398__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__397__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__396__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_165_)
);

scs8hd_diode_2 ANTENNA__408__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__407__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__406__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__405__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__404__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__403__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_166_)
);

scs8hd_diode_2 ANTENNA__415__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__414__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__413__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__412__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__411__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__410__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_167_)
);

scs8hd_diode_2 ANTENNA__422__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__421__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__420__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__419__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__418__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__417__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_168_)
);

scs8hd_diode_2 ANTENNA__433__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_169_)
);

scs8hd_diode_2 ANTENNA__432__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_169_)
);

scs8hd_diode_2 ANTENNA__433__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_170_)
);

scs8hd_diode_2 ANTENNA__432__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_170_)
);

scs8hd_diode_2 ANTENNA__561__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__518__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__475__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__435__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__429__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__345__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_171_)
);

scs8hd_diode_2 ANTENNA__468__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__461__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__454__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__447__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__440__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__430__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_172_)
);

scs8hd_diode_2 ANTENNA__431__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_173_)
);

scs8hd_diode_2 ANTENNA__434__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_174_)
);

scs8hd_diode_2 ANTENNA__433__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_174_)
);

scs8hd_diode_2 ANTENNA__434__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_175_)
);

scs8hd_diode_2 ANTENNA__433__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_175_)
);

scs8hd_diode_2 ANTENNA__437__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_176_)
);

scs8hd_diode_2 ANTENNA__436__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_176_)
);

scs8hd_diode_2 ANTENNA__443__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_177_)
);

scs8hd_diode_2 ANTENNA__442__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_177_)
);

scs8hd_diode_2 ANTENNA__443__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_178_)
);

scs8hd_diode_2 ANTENNA__442__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_178_)
);

scs8hd_diode_2 ANTENNA__441__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_179_)
);

scs8hd_diode_2 ANTENNA__444__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_180_)
);

scs8hd_diode_2 ANTENNA__443__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_180_)
);

scs8hd_diode_2 ANTENNA__444__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_181_)
);

scs8hd_diode_2 ANTENNA__443__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_181_)
);

scs8hd_diode_2 ANTENNA__450__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_182_)
);

scs8hd_diode_2 ANTENNA__449__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_182_)
);

scs8hd_diode_2 ANTENNA__450__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_183_)
);

scs8hd_diode_2 ANTENNA__449__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_183_)
);

scs8hd_diode_2 ANTENNA__448__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_184_)
);

scs8hd_diode_2 ANTENNA__451__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_185_)
);

scs8hd_diode_2 ANTENNA__450__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_185_)
);

scs8hd_diode_2 ANTENNA__451__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_186_)
);

scs8hd_diode_2 ANTENNA__450__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_186_)
);

scs8hd_diode_2 ANTENNA__457__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_187_)
);

scs8hd_diode_2 ANTENNA__456__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_187_)
);

scs8hd_diode_2 ANTENNA__457__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_188_)
);

scs8hd_diode_2 ANTENNA__456__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_188_)
);

scs8hd_diode_2 ANTENNA__455__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_189_)
);

scs8hd_diode_2 ANTENNA__458__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_190_)
);

scs8hd_diode_2 ANTENNA__457__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_190_)
);

scs8hd_diode_2 ANTENNA__458__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_191_)
);

scs8hd_diode_2 ANTENNA__457__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_191_)
);

scs8hd_diode_2 ANTENNA__464__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_192_)
);

scs8hd_diode_2 ANTENNA__463__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_192_)
);

scs8hd_diode_2 ANTENNA__464__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_193_)
);

scs8hd_diode_2 ANTENNA__463__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_193_)
);

scs8hd_diode_2 ANTENNA__462__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_194_)
);

scs8hd_diode_2 ANTENNA__465__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_195_)
);

scs8hd_diode_2 ANTENNA__464__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_195_)
);

scs8hd_diode_2 ANTENNA__465__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_196_)
);

scs8hd_diode_2 ANTENNA__464__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_196_)
);

scs8hd_diode_2 ANTENNA__471__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_197_)
);

scs8hd_diode_2 ANTENNA__470__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_197_)
);

scs8hd_diode_2 ANTENNA__471__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_198_)
);

scs8hd_diode_2 ANTENNA__470__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_198_)
);

scs8hd_diode_2 ANTENNA__469__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_199_)
);

scs8hd_diode_2 ANTENNA__472__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_200_)
);

scs8hd_diode_2 ANTENNA__471__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_200_)
);

scs8hd_diode_2 ANTENNA__472__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_201_)
);

scs8hd_diode_2 ANTENNA__471__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_201_)
);

scs8hd_diode_2 ANTENNA__479__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_202_)
);

scs8hd_diode_2 ANTENNA__478__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_202_)
);

scs8hd_diode_2 ANTENNA__479__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_203_)
);

scs8hd_diode_2 ANTENNA__478__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_203_)
);

scs8hd_diode_2 ANTENNA__511__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__504__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__497__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__490__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__483__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__476__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_204_)
);

scs8hd_diode_2 ANTENNA__477__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_205_)
);

scs8hd_diode_2 ANTENNA__480__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_206_)
);

scs8hd_diode_2 ANTENNA__479__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_206_)
);

scs8hd_diode_2 ANTENNA__480__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_207_)
);

scs8hd_diode_2 ANTENNA__479__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_207_)
);

scs8hd_diode_2 ANTENNA__486__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_208_)
);

scs8hd_diode_2 ANTENNA__485__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_208_)
);

scs8hd_diode_2 ANTENNA__486__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_209_)
);

scs8hd_diode_2 ANTENNA__485__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_209_)
);

scs8hd_diode_2 ANTENNA__484__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_210_)
);

scs8hd_diode_2 ANTENNA__487__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_211_)
);

scs8hd_diode_2 ANTENNA__486__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_211_)
);

scs8hd_diode_2 ANTENNA__487__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_212_)
);

scs8hd_diode_2 ANTENNA__486__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_212_)
);

scs8hd_diode_2 ANTENNA__493__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_213_)
);

scs8hd_diode_2 ANTENNA__492__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_213_)
);

scs8hd_diode_2 ANTENNA__493__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_214_)
);

scs8hd_diode_2 ANTENNA__492__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_214_)
);

scs8hd_diode_2 ANTENNA__491__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_215_)
);

scs8hd_diode_2 ANTENNA__494__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_216_)
);

scs8hd_diode_2 ANTENNA__493__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_216_)
);

scs8hd_diode_2 ANTENNA__494__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_217_)
);

scs8hd_diode_2 ANTENNA__493__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_217_)
);

scs8hd_diode_2 ANTENNA__500__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_218_)
);

scs8hd_diode_2 ANTENNA__499__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_218_)
);

scs8hd_diode_2 ANTENNA__500__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_219_)
);

scs8hd_diode_2 ANTENNA__499__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_219_)
);

scs8hd_diode_2 ANTENNA__498__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_220_)
);

scs8hd_diode_2 ANTENNA__501__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_221_)
);

scs8hd_diode_2 ANTENNA__500__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_221_)
);

scs8hd_diode_2 ANTENNA__501__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_222_)
);

scs8hd_diode_2 ANTENNA__500__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_222_)
);

scs8hd_diode_2 ANTENNA__507__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_223_)
);

scs8hd_diode_2 ANTENNA__506__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_223_)
);

scs8hd_diode_2 ANTENNA__507__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_224_)
);

scs8hd_diode_2 ANTENNA__506__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_224_)
);

scs8hd_diode_2 ANTENNA__505__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_225_)
);

scs8hd_diode_2 ANTENNA__508__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_226_)
);

scs8hd_diode_2 ANTENNA__507__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_226_)
);

scs8hd_diode_2 ANTENNA__508__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_227_)
);

scs8hd_diode_2 ANTENNA__507__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_227_)
);

scs8hd_diode_2 ANTENNA__514__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_228_)
);

scs8hd_diode_2 ANTENNA__513__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_228_)
);

scs8hd_diode_2 ANTENNA__514__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_229_)
);

scs8hd_diode_2 ANTENNA__513__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_229_)
);

scs8hd_diode_2 ANTENNA__512__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_230_)
);

scs8hd_diode_2 ANTENNA__515__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_231_)
);

scs8hd_diode_2 ANTENNA__514__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_231_)
);

scs8hd_diode_2 ANTENNA__515__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_232_)
);

scs8hd_diode_2 ANTENNA__514__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_232_)
);

scs8hd_diode_2 ANTENNA__522__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_233_)
);

scs8hd_diode_2 ANTENNA__521__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_233_)
);

scs8hd_diode_2 ANTENNA__522__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_234_)
);

scs8hd_diode_2 ANTENNA__521__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_234_)
);

scs8hd_diode_2 ANTENNA__554__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__547__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__540__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__533__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__526__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__519__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_235_)
);

scs8hd_diode_2 ANTENNA__520__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_236_)
);

scs8hd_diode_2 ANTENNA__523__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_237_)
);

scs8hd_diode_2 ANTENNA__522__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_237_)
);

scs8hd_diode_2 ANTENNA__523__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_238_)
);

scs8hd_diode_2 ANTENNA__522__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_238_)
);

scs8hd_diode_2 ANTENNA__529__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_239_)
);

scs8hd_diode_2 ANTENNA__528__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_239_)
);

scs8hd_diode_2 ANTENNA__529__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_240_)
);

scs8hd_diode_2 ANTENNA__528__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_240_)
);

scs8hd_diode_2 ANTENNA__527__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_241_)
);

scs8hd_diode_2 ANTENNA__530__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_242_)
);

scs8hd_diode_2 ANTENNA__529__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_242_)
);

scs8hd_diode_2 ANTENNA__530__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_243_)
);

scs8hd_diode_2 ANTENNA__529__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_243_)
);

scs8hd_diode_2 ANTENNA__536__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_244_)
);

scs8hd_diode_2 ANTENNA__535__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_244_)
);

scs8hd_diode_2 ANTENNA__536__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_245_)
);

scs8hd_diode_2 ANTENNA__535__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_245_)
);

scs8hd_diode_2 ANTENNA__534__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_246_)
);

scs8hd_diode_2 ANTENNA__537__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_247_)
);

scs8hd_diode_2 ANTENNA__536__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_247_)
);

scs8hd_diode_2 ANTENNA__537__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_248_)
);

scs8hd_diode_2 ANTENNA__536__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_248_)
);

scs8hd_diode_2 ANTENNA__543__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_249_)
);

scs8hd_diode_2 ANTENNA__542__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_249_)
);

scs8hd_diode_2 ANTENNA__543__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_250_)
);

scs8hd_diode_2 ANTENNA__542__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_250_)
);

scs8hd_diode_2 ANTENNA__541__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_251_)
);

scs8hd_diode_2 ANTENNA__544__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_252_)
);

scs8hd_diode_2 ANTENNA__543__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_252_)
);

scs8hd_diode_2 ANTENNA__544__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_253_)
);

scs8hd_diode_2 ANTENNA__543__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_253_)
);

scs8hd_diode_2 ANTENNA__550__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_254_)
);

scs8hd_diode_2 ANTENNA__549__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_254_)
);

scs8hd_diode_2 ANTENNA__550__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_255_)
);

scs8hd_diode_2 ANTENNA__549__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_255_)
);

scs8hd_diode_2 ANTENNA__548__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_256_)
);

scs8hd_diode_2 ANTENNA__551__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_257_)
);

scs8hd_diode_2 ANTENNA__550__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_257_)
);

scs8hd_diode_2 ANTENNA__551__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_258_)
);

scs8hd_diode_2 ANTENNA__550__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_258_)
);

scs8hd_diode_2 ANTENNA__557__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_259_)
);

scs8hd_diode_2 ANTENNA__556__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_259_)
);

scs8hd_diode_2 ANTENNA__557__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_260_)
);

scs8hd_diode_2 ANTENNA__556__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_260_)
);

scs8hd_diode_2 ANTENNA__555__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_261_)
);

scs8hd_diode_2 ANTENNA__558__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_262_)
);

scs8hd_diode_2 ANTENNA__557__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_262_)
);

scs8hd_diode_2 ANTENNA__558__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_263_)
);

scs8hd_diode_2 ANTENNA__557__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_263_)
);

scs8hd_diode_2 ANTENNA__565__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_264_)
);

scs8hd_diode_2 ANTENNA__564__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_264_)
);

scs8hd_diode_2 ANTENNA__565__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_265_)
);

scs8hd_diode_2 ANTENNA__564__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_265_)
);

scs8hd_diode_2 ANTENNA__597__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__590__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__583__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__576__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__569__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__562__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_266_)
);

scs8hd_diode_2 ANTENNA__563__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_267_)
);

scs8hd_diode_2 ANTENNA__566__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_268_)
);

scs8hd_diode_2 ANTENNA__565__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_268_)
);

scs8hd_diode_2 ANTENNA__566__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_269_)
);

scs8hd_diode_2 ANTENNA__565__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_269_)
);

scs8hd_diode_2 ANTENNA__572__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_270_)
);

scs8hd_diode_2 ANTENNA__571__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_270_)
);

scs8hd_diode_2 ANTENNA__572__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_271_)
);

scs8hd_diode_2 ANTENNA__571__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_271_)
);

scs8hd_diode_2 ANTENNA__570__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_272_)
);

scs8hd_diode_2 ANTENNA__573__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_273_)
);

scs8hd_diode_2 ANTENNA__572__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_273_)
);

scs8hd_diode_2 ANTENNA__573__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_274_)
);

scs8hd_diode_2 ANTENNA__572__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_274_)
);

scs8hd_diode_2 ANTENNA__579__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_275_)
);

scs8hd_diode_2 ANTENNA__578__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_275_)
);

scs8hd_diode_2 ANTENNA__579__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_276_)
);

scs8hd_diode_2 ANTENNA__578__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_276_)
);

scs8hd_diode_2 ANTENNA__577__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_277_)
);

scs8hd_diode_2 ANTENNA__580__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_278_)
);

scs8hd_diode_2 ANTENNA__579__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_278_)
);

scs8hd_diode_2 ANTENNA__580__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_279_)
);

scs8hd_diode_2 ANTENNA__579__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_279_)
);

scs8hd_diode_2 ANTENNA__586__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_280_)
);

scs8hd_diode_2 ANTENNA__585__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_280_)
);

scs8hd_diode_2 ANTENNA__586__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_281_)
);

scs8hd_diode_2 ANTENNA__585__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_281_)
);

scs8hd_diode_2 ANTENNA__584__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_282_)
);

scs8hd_diode_2 ANTENNA__587__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_283_)
);

scs8hd_diode_2 ANTENNA__586__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_283_)
);

scs8hd_diode_2 ANTENNA__587__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_284_)
);

scs8hd_diode_2 ANTENNA__586__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_284_)
);

scs8hd_diode_2 ANTENNA__593__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_285_)
);

scs8hd_diode_2 ANTENNA__592__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_285_)
);

scs8hd_diode_2 ANTENNA__593__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_286_)
);

scs8hd_diode_2 ANTENNA__592__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_286_)
);

scs8hd_diode_2 ANTENNA__591__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_287_)
);

scs8hd_diode_2 ANTENNA__594__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_288_)
);

scs8hd_diode_2 ANTENNA__593__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_288_)
);

scs8hd_diode_2 ANTENNA__594__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_289_)
);

scs8hd_diode_2 ANTENNA__593__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_289_)
);

scs8hd_diode_2 ANTENNA__600__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_290_)
);

scs8hd_diode_2 ANTENNA__599__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_290_)
);

scs8hd_diode_2 ANTENNA__600__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_291_)
);

scs8hd_diode_2 ANTENNA__599__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_291_)
);

scs8hd_diode_2 ANTENNA__598__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_292_)
);

scs8hd_diode_2 ANTENNA__601__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_293_)
);

scs8hd_diode_2 ANTENNA__600__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_293_)
);

scs8hd_diode_2 ANTENNA__601__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_294_)
);

scs8hd_diode_2 ANTENNA__600__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_294_)
);

scs8hd_diode_2 ANTENNA__608__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_295_)
);

scs8hd_diode_2 ANTENNA__607__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_295_)
);

scs8hd_diode_2 ANTENNA__608__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_296_)
);

scs8hd_diode_2 ANTENNA__607__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_296_)
);

scs8hd_diode_2 ANTENNA__626__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__619__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__612__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__605__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__338__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__331__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_297_)
);

scs8hd_diode_2 ANTENNA__606__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_298_)
);

scs8hd_diode_2 ANTENNA__609__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_299_)
);

scs8hd_diode_2 ANTENNA__608__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_299_)
);

scs8hd_diode_2 ANTENNA__609__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_300_)
);

scs8hd_diode_2 ANTENNA__608__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_300_)
);

scs8hd_diode_2 ANTENNA__615__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_301_)
);

scs8hd_diode_2 ANTENNA__614__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_301_)
);

scs8hd_diode_2 ANTENNA__615__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_302_)
);

scs8hd_diode_2 ANTENNA__614__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_302_)
);

scs8hd_diode_2 ANTENNA__613__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_303_)
);

scs8hd_diode_2 ANTENNA__616__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_304_)
);

scs8hd_diode_2 ANTENNA__615__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_304_)
);

scs8hd_diode_2 ANTENNA__616__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_305_)
);

scs8hd_diode_2 ANTENNA__615__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_305_)
);

scs8hd_diode_2 ANTENNA__622__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_306_)
);

scs8hd_diode_2 ANTENNA__621__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_306_)
);

scs8hd_diode_2 ANTENNA__622__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_307_)
);

scs8hd_diode_2 ANTENNA__621__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_307_)
);

scs8hd_diode_2 ANTENNA__620__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_308_)
);

scs8hd_diode_2 ANTENNA__623__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_309_)
);

scs8hd_diode_2 ANTENNA__622__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_309_)
);

scs8hd_diode_2 ANTENNA__623__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_310_)
);

scs8hd_diode_2 ANTENNA__622__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_310_)
);

scs8hd_diode_2 ANTENNA__629__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_311_)
);

scs8hd_diode_2 ANTENNA__628__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_311_)
);

scs8hd_diode_2 ANTENNA__629__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_312_)
);

scs8hd_diode_2 ANTENNA__628__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_312_)
);

scs8hd_diode_2 ANTENNA__627__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_313_)
);

scs8hd_diode_2 ANTENNA__630__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_314_)
);

scs8hd_diode_2 ANTENNA__629__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_314_)
);

scs8hd_diode_2 ANTENNA__630__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_315_)
);

scs8hd_diode_2 ANTENNA__629__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_315_)
);

scs8hd_diode_2 ANTENNA__334__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_316_)
);

scs8hd_diode_2 ANTENNA__333__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_316_)
);

scs8hd_diode_2 ANTENNA__334__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_317_)
);

scs8hd_diode_2 ANTENNA__333__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_317_)
);

scs8hd_diode_2 ANTENNA__332__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_318_)
);

scs8hd_diode_2 ANTENNA__335__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_319_)
);

scs8hd_diode_2 ANTENNA__334__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_319_)
);

scs8hd_diode_2 ANTENNA__335__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_320_)
);

scs8hd_diode_2 ANTENNA__334__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_320_)
);

scs8hd_diode_2 ANTENNA__341__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_321_)
);

scs8hd_diode_2 ANTENNA__340__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_321_)
);

scs8hd_diode_2 ANTENNA__341__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_322_)
);

scs8hd_diode_2 ANTENNA__340__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_322_)
);

scs8hd_diode_2 ANTENNA__339__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_323_)
);

scs8hd_diode_2 ANTENNA__342__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_324_)
);

scs8hd_diode_2 ANTENNA__341__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_324_)
);

scs8hd_diode_2 ANTENNA__342__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_325_)
);

scs8hd_diode_2 ANTENNA__341__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_325_)
);

scs8hd_diode_2 ANTENNA__348__A1N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_326_)
);

scs8hd_diode_2 ANTENNA__347__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_326_)
);

scs8hd_diode_2 ANTENNA__348__A2N (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_327_)
);

scs8hd_diode_2 ANTENNA__347__A2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_327_)
);

scs8hd_diode_2 ANTENNA__346__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_328_)
);

scs8hd_diode_2 ANTENNA__349__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_329_)
);

scs8hd_diode_2 ANTENNA__348__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_329_)
);

scs8hd_diode_2 ANTENNA__349__B (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_330_)
);

scs8hd_diode_2 ANTENNA__348__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(_330_)
);

scs8hd_diode_2 ANTENNA__648__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__647__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__646__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__645__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__644__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__643__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__642__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__641__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__640__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__639__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__638__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__637__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__636__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__635__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__634__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__633__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_0)
);

scs8hd_diode_2 ANTENNA__664__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__663__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__662__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__661__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__660__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__659__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__658__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__657__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__656__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__655__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__654__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__653__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__652__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__651__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__650__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__649__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_16)
);

scs8hd_diode_2 ANTENNA__680__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__679__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__678__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__677__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__676__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__675__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__674__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__673__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__672__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__671__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__670__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__669__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__668__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__667__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__666__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__665__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_32)
);

scs8hd_diode_2 ANTENNA__696__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__695__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__694__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__693__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__692__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__691__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__690__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__689__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__688__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__687__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__686__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__685__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__684__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__683__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__682__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__681__CLK (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_0_48)
);

scs8hd_diode_2 ANTENNA__CTS_buf_1_48_A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_1_0)
);

scs8hd_diode_2 ANTENNA__CTS_buf_1_32_A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_1_0)
);

scs8hd_diode_2 ANTENNA__CTS_buf_1_16_A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_1_0)
);

scs8hd_diode_2 ANTENNA__CTS_buf_1_0_A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(clk_1_0)
);

scs8hd_diode_2 ANTENNA__634__D (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\csa0.hsum2 )
);

scs8hd_diode_2 ANTENNA__432__B1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\csa0.sc )
);

scs8hd_diode_2 ANTENNA__426__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\csa0.sc )
);

scs8hd_diode_2 ANTENNA__432__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\csa0.y )
);

scs8hd_diode_2 ANTENNA__427__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\csa0.y )
);

scs8hd_diode_2 ANTENNA__499__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[10] )
);

scs8hd_diode_2 ANTENNA__496__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[10] )
);

scs8hd_diode_2 ANTENNA__506__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[11] )
);

scs8hd_diode_2 ANTENNA__503__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[11] )
);

scs8hd_diode_2 ANTENNA__513__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[12] )
);

scs8hd_diode_2 ANTENNA__510__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[12] )
);

scs8hd_diode_2 ANTENNA__521__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[13] )
);

scs8hd_diode_2 ANTENNA__517__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[13] )
);

scs8hd_diode_2 ANTENNA__528__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[14] )
);

scs8hd_diode_2 ANTENNA__525__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[14] )
);

scs8hd_diode_2 ANTENNA__535__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[15] )
);

scs8hd_diode_2 ANTENNA__532__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[15] )
);

scs8hd_diode_2 ANTENNA__542__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[16] )
);

scs8hd_diode_2 ANTENNA__539__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[16] )
);

scs8hd_diode_2 ANTENNA__549__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[17] )
);

scs8hd_diode_2 ANTENNA__546__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[17] )
);

scs8hd_diode_2 ANTENNA__556__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[18] )
);

scs8hd_diode_2 ANTENNA__553__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[18] )
);

scs8hd_diode_2 ANTENNA__564__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[19] )
);

scs8hd_diode_2 ANTENNA__560__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[19] )
);

scs8hd_diode_2 ANTENNA__571__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[20] )
);

scs8hd_diode_2 ANTENNA__568__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[20] )
);

scs8hd_diode_2 ANTENNA__578__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[21] )
);

scs8hd_diode_2 ANTENNA__575__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[21] )
);

scs8hd_diode_2 ANTENNA__585__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[22] )
);

scs8hd_diode_2 ANTENNA__582__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[22] )
);

scs8hd_diode_2 ANTENNA__592__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[23] )
);

scs8hd_diode_2 ANTENNA__589__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[23] )
);

scs8hd_diode_2 ANTENNA__599__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[24] )
);

scs8hd_diode_2 ANTENNA__596__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[24] )
);

scs8hd_diode_2 ANTENNA__607__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[25] )
);

scs8hd_diode_2 ANTENNA__603__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[25] )
);

scs8hd_diode_2 ANTENNA__614__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[26] )
);

scs8hd_diode_2 ANTENNA__611__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[26] )
);

scs8hd_diode_2 ANTENNA__621__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[27] )
);

scs8hd_diode_2 ANTENNA__618__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[27] )
);

scs8hd_diode_2 ANTENNA__628__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[28] )
);

scs8hd_diode_2 ANTENNA__625__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[28] )
);

scs8hd_diode_2 ANTENNA__632__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[29] )
);

scs8hd_diode_2 ANTENNA__333__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[29] )
);

scs8hd_diode_2 ANTENNA__442__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[2] )
);

scs8hd_diode_2 ANTENNA__439__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[2] )
);

scs8hd_diode_2 ANTENNA__340__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[30] )
);

scs8hd_diode_2 ANTENNA__337__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[30] )
);

scs8hd_diode_2 ANTENNA__449__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[3] )
);

scs8hd_diode_2 ANTENNA__446__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[3] )
);

scs8hd_diode_2 ANTENNA__456__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[4] )
);

scs8hd_diode_2 ANTENNA__453__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[4] )
);

scs8hd_diode_2 ANTENNA__463__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[5] )
);

scs8hd_diode_2 ANTENNA__460__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[5] )
);

scs8hd_diode_2 ANTENNA__470__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[6] )
);

scs8hd_diode_2 ANTENNA__467__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[6] )
);

scs8hd_diode_2 ANTENNA__478__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[7] )
);

scs8hd_diode_2 ANTENNA__474__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[7] )
);

scs8hd_diode_2 ANTENNA__485__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[8] )
);

scs8hd_diode_2 ANTENNA__482__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[8] )
);

scs8hd_diode_2 ANTENNA__492__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[9] )
);

scs8hd_diode_2 ANTENNA__489__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\pp[9] )
);

scs8hd_diode_2 ANTENNA__347__B2 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\tcmp.s )
);

scs8hd_diode_2 ANTENNA__344__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\tcmp.s )
);

scs8hd_diode_2 ANTENNA__437__A1 (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\tcmp.z )
);

scs8hd_diode_2 ANTENNA__436__A (
    .vpwr(vpwr),
    .vgnd(vgnd),
    .DIODE(\tcmp.z )
);

endmodule
