magic
tech EFS8A
magscale 1 2
timestamp 1595162803
<< locali >>
rect 13185 22627 13219 22661
rect 13185 22593 13311 22627
rect 16589 16031 16623 16201
rect 13185 14535 13219 14569
rect 13093 14501 13219 14535
rect 4077 14399 4111 14501
rect 3433 12631 3467 12869
rect 9505 11679 9539 11781
rect 10241 11611 10275 11713
rect 4169 2499 4203 2601
rect 4169 2465 4287 2499
<< viali >>
rect 4997 25313 5031 25347
rect 8401 25313 8435 25347
rect 12265 25313 12299 25347
rect 13093 25313 13127 25347
rect 15669 25313 15703 25347
rect 16773 25313 16807 25347
rect 22385 25313 22419 25347
rect 22845 25313 22879 25347
rect 4905 25245 4939 25279
rect 5733 25245 5767 25279
rect 8309 25245 8343 25279
rect 14105 25177 14139 25211
rect 15853 25177 15887 25211
rect 5181 25109 5215 25143
rect 8585 25109 8619 25143
rect 10057 25109 10091 25143
rect 10885 25109 10919 25143
rect 13461 25109 13495 25143
rect 14473 25109 14507 25143
rect 16957 25109 16991 25143
rect 22569 25109 22603 25143
rect 4905 24905 4939 24939
rect 7297 24905 7331 24939
rect 8309 24905 8343 24939
rect 16129 24905 16163 24939
rect 16773 24905 16807 24939
rect 22477 24905 22511 24939
rect 23121 24905 23155 24939
rect 7757 24769 7791 24803
rect 9413 24769 9447 24803
rect 12633 24769 12667 24803
rect 13185 24769 13219 24803
rect 3893 24701 3927 24735
rect 4169 24701 4203 24735
rect 5825 24701 5859 24735
rect 6193 24701 6227 24735
rect 8033 24701 8067 24735
rect 8125 24701 8159 24735
rect 9505 24701 9539 24735
rect 10333 24701 10367 24735
rect 10885 24701 10919 24735
rect 12725 24701 12759 24735
rect 13461 24701 13495 24735
rect 14197 24701 14231 24735
rect 14565 24701 14599 24735
rect 18889 24701 18923 24735
rect 19625 24701 19659 24735
rect 20913 24701 20947 24735
rect 21189 24701 21223 24735
rect 22201 24701 22235 24735
rect 22293 24701 22327 24735
rect 9965 24633 9999 24667
rect 11529 24633 11563 24667
rect 12081 24633 12115 24667
rect 17693 24633 17727 24667
rect 4353 24565 4387 24599
rect 5457 24565 5491 24599
rect 8953 24565 8987 24599
rect 17325 24565 17359 24599
rect 21373 24565 21407 24599
rect 21833 24565 21867 24599
rect 9045 24361 9079 24395
rect 14841 24361 14875 24395
rect 17877 24361 17911 24395
rect 15761 24293 15795 24327
rect 17233 24293 17267 24327
rect 1685 24225 1719 24259
rect 4629 24225 4663 24259
rect 4721 24225 4755 24259
rect 5181 24225 5215 24259
rect 5365 24225 5399 24259
rect 6377 24225 6411 24259
rect 6745 24225 6779 24259
rect 7665 24225 7699 24259
rect 8309 24225 8343 24259
rect 10977 24225 11011 24259
rect 11437 24225 11471 24259
rect 12955 24225 12989 24259
rect 13461 24225 13495 24259
rect 13553 24225 13587 24259
rect 14565 24225 14599 24259
rect 16405 24225 16439 24259
rect 16773 24225 16807 24259
rect 16957 24225 16991 24259
rect 18797 24225 18831 24259
rect 18889 24225 18923 24259
rect 19349 24225 19383 24259
rect 19533 24225 19567 24259
rect 21189 24225 21223 24259
rect 22661 24225 22695 24259
rect 1593 24157 1627 24191
rect 7389 24157 7423 24191
rect 8217 24157 8251 24191
rect 8769 24157 8803 24191
rect 12817 24157 12851 24191
rect 16497 24157 16531 24191
rect 18337 24157 18371 24191
rect 21097 24157 21131 24191
rect 22569 24157 22603 24191
rect 5549 24089 5583 24123
rect 13921 24089 13955 24123
rect 19717 24089 19751 24123
rect 1869 24021 1903 24055
rect 2605 24021 2639 24055
rect 11989 24021 12023 24055
rect 12449 24021 12483 24055
rect 22845 24021 22879 24055
rect 1685 23817 1719 23851
rect 2053 23817 2087 23851
rect 4813 23817 4847 23851
rect 6377 23817 6411 23851
rect 8493 23817 8527 23851
rect 8953 23817 8987 23851
rect 9781 23817 9815 23851
rect 10517 23817 10551 23851
rect 11713 23817 11747 23851
rect 15209 23817 15243 23851
rect 17509 23817 17543 23851
rect 18889 23817 18923 23851
rect 20913 23817 20947 23851
rect 22661 23817 22695 23851
rect 22937 23817 22971 23851
rect 5457 23749 5491 23783
rect 10885 23749 10919 23783
rect 11345 23749 11379 23783
rect 17141 23749 17175 23783
rect 5181 23681 5215 23715
rect 6101 23681 6135 23715
rect 12081 23681 12115 23715
rect 12909 23681 12943 23715
rect 15485 23681 15519 23715
rect 19165 23681 19199 23715
rect 19717 23681 19751 23715
rect 2973 23613 3007 23647
rect 3157 23613 3191 23647
rect 7481 23613 7515 23647
rect 7665 23613 7699 23647
rect 7987 23613 8021 23647
rect 8125 23613 8159 23647
rect 9597 23613 9631 23647
rect 10057 23613 10091 23647
rect 12633 23613 12667 23647
rect 15669 23613 15703 23647
rect 16129 23613 16163 23647
rect 16221 23613 16255 23647
rect 19809 23613 19843 23647
rect 20177 23613 20211 23647
rect 20361 23613 20395 23647
rect 21833 23613 21867 23647
rect 22201 23613 22235 23647
rect 7021 23545 7055 23579
rect 14657 23545 14691 23579
rect 18521 23545 18555 23579
rect 21189 23545 21223 23579
rect 16681 23477 16715 23511
rect 2605 23273 2639 23307
rect 4445 23273 4479 23307
rect 7113 23273 7147 23307
rect 11621 23273 11655 23307
rect 12265 23273 12299 23307
rect 13829 23273 13863 23307
rect 15577 23273 15611 23307
rect 18521 23273 18555 23307
rect 19165 23273 19199 23307
rect 19993 23273 20027 23307
rect 4997 23205 5031 23239
rect 6745 23205 6779 23239
rect 18889 23205 18923 23239
rect 19625 23205 19659 23239
rect 1593 23137 1627 23171
rect 7573 23137 7607 23171
rect 8585 23137 8619 23171
rect 9321 23137 9355 23171
rect 9873 23137 9907 23171
rect 12633 23137 12667 23171
rect 13001 23137 13035 23171
rect 23029 23137 23063 23171
rect 2237 23069 2271 23103
rect 4721 23069 4755 23103
rect 12449 23069 12483 23103
rect 12909 23069 12943 23103
rect 13461 23069 13495 23103
rect 14289 23069 14323 23103
rect 15945 23069 15979 23103
rect 16221 23069 16255 23103
rect 17969 23069 18003 23103
rect 21465 23069 21499 23103
rect 22845 23069 22879 23103
rect 10793 23001 10827 23035
rect 22109 23001 22143 23035
rect 1777 22933 1811 22967
rect 2973 22933 3007 22967
rect 7757 22933 7791 22967
rect 8769 22933 8803 22967
rect 10057 22933 10091 22967
rect 10425 22933 10459 22967
rect 11069 22933 11103 22967
rect 14933 22933 14967 22967
rect 21741 22933 21775 22967
rect 4813 22729 4847 22763
rect 5181 22729 5215 22763
rect 5733 22729 5767 22763
rect 7205 22729 7239 22763
rect 11989 22729 12023 22763
rect 15853 22729 15887 22763
rect 23029 22729 23063 22763
rect 13185 22661 13219 22695
rect 1869 22593 1903 22627
rect 2421 22593 2455 22627
rect 9965 22593 9999 22627
rect 10701 22593 10735 22627
rect 11161 22593 11195 22627
rect 16129 22593 16163 22627
rect 18705 22593 18739 22627
rect 20453 22593 20487 22627
rect 2145 22525 2179 22559
rect 5549 22525 5583 22559
rect 7941 22525 7975 22559
rect 8401 22525 8435 22559
rect 10885 22525 10919 22559
rect 11253 22525 11287 22559
rect 16313 22525 16347 22559
rect 17325 22525 17359 22559
rect 18429 22525 18463 22559
rect 21373 22525 21407 22559
rect 21557 22525 21591 22559
rect 22109 22525 22143 22559
rect 22293 22525 22327 22559
rect 4169 22457 4203 22491
rect 10241 22457 10275 22491
rect 13001 22457 13035 22491
rect 13553 22457 13587 22491
rect 15301 22457 15335 22491
rect 21097 22457 21131 22491
rect 6009 22389 6043 22423
rect 6377 22389 6411 22423
rect 17693 22389 17727 22423
rect 22569 22389 22603 22423
rect 1593 22185 1627 22219
rect 3525 22185 3559 22219
rect 4261 22185 4295 22219
rect 7573 22185 7607 22219
rect 8585 22185 8619 22219
rect 11621 22185 11655 22219
rect 13369 22185 13403 22219
rect 14381 22185 14415 22219
rect 14749 22185 14783 22219
rect 16037 22185 16071 22219
rect 16773 22185 16807 22219
rect 9321 22117 9355 22151
rect 11897 22117 11931 22151
rect 19901 22117 19935 22151
rect 20545 22117 20579 22151
rect 3065 22049 3099 22083
rect 5365 22049 5399 22083
rect 6101 22049 6135 22083
rect 7941 22049 7975 22083
rect 10057 22049 10091 22083
rect 10517 22049 10551 22083
rect 10609 22049 10643 22083
rect 12541 22049 12575 22083
rect 14197 22049 14231 22083
rect 16589 22049 16623 22083
rect 17601 22049 17635 22083
rect 17877 22049 17911 22083
rect 21189 22049 21223 22083
rect 21741 22049 21775 22083
rect 2421 21981 2455 22015
rect 9965 21981 9999 22015
rect 12909 21981 12943 22015
rect 13737 21981 13771 22015
rect 15669 21981 15703 22015
rect 18153 21981 18187 22015
rect 10977 21913 11011 21947
rect 2053 21845 2087 21879
rect 23305 21845 23339 21879
rect 4169 21641 4203 21675
rect 5273 21641 5307 21675
rect 8401 21641 8435 21675
rect 11989 21641 12023 21675
rect 16221 21641 16255 21675
rect 17693 21641 17727 21675
rect 23029 21641 23063 21675
rect 4905 21573 4939 21607
rect 17325 21573 17359 21607
rect 20269 21573 20303 21607
rect 21281 21573 21315 21607
rect 2881 21505 2915 21539
rect 9137 21505 9171 21539
rect 9689 21505 9723 21539
rect 11437 21505 11471 21539
rect 12909 21505 12943 21539
rect 14657 21505 14691 21539
rect 19165 21505 19199 21539
rect 21557 21505 21591 21539
rect 22293 21505 22327 21539
rect 1685 21437 1719 21471
rect 2421 21437 2455 21471
rect 2605 21437 2639 21471
rect 2973 21437 3007 21471
rect 3985 21437 4019 21471
rect 9413 21437 9447 21471
rect 12633 21437 12667 21471
rect 18705 21437 18739 21471
rect 18889 21437 18923 21471
rect 19257 21437 19291 21471
rect 20085 21437 20119 21471
rect 22201 21437 22235 21471
rect 22569 21437 22603 21471
rect 22753 21437 22787 21471
rect 3433 21369 3467 21403
rect 8769 21369 8803 21403
rect 18245 21369 18279 21403
rect 19717 21369 19751 21403
rect 2237 21301 2271 21335
rect 4537 21301 4571 21335
rect 14933 21301 14967 21335
rect 16589 21301 16623 21335
rect 20637 21301 20671 21335
rect 3617 21097 3651 21131
rect 8585 21097 8619 21131
rect 8861 21097 8895 21131
rect 12357 21097 12391 21131
rect 12725 21097 12759 21131
rect 13369 21097 13403 21131
rect 14749 21097 14783 21131
rect 18337 21097 18371 21131
rect 20545 21097 20579 21131
rect 21281 21097 21315 21131
rect 3249 21029 3283 21063
rect 5641 21029 5675 21063
rect 7389 21029 7423 21063
rect 9321 21029 9355 21063
rect 9965 21029 9999 21063
rect 11897 21029 11931 21063
rect 17969 21029 18003 21063
rect 21833 21029 21867 21063
rect 1777 20961 1811 20995
rect 2329 20961 2363 20995
rect 2513 20961 2547 20995
rect 4261 20961 4295 20995
rect 10425 20961 10459 20995
rect 12173 20961 12207 20995
rect 13185 20961 13219 20995
rect 14197 20961 14231 20995
rect 16497 20961 16531 20995
rect 16957 20961 16991 20995
rect 19625 20961 19659 20995
rect 1685 20893 1719 20927
rect 5365 20893 5399 20927
rect 18981 20893 19015 20927
rect 20085 20893 20119 20927
rect 21557 20893 21591 20927
rect 23581 20893 23615 20927
rect 2697 20825 2731 20859
rect 4445 20825 4479 20859
rect 7941 20825 7975 20859
rect 14381 20825 14415 20859
rect 18613 20757 18647 20791
rect 5457 20553 5491 20587
rect 10885 20553 10919 20587
rect 16405 20553 16439 20587
rect 16773 20553 16807 20587
rect 17049 20553 17083 20587
rect 18337 20553 18371 20587
rect 21925 20553 21959 20587
rect 22385 20553 22419 20587
rect 10241 20485 10275 20519
rect 1869 20417 1903 20451
rect 2421 20417 2455 20451
rect 4169 20417 4203 20451
rect 7573 20417 7607 20451
rect 8125 20417 8159 20451
rect 14013 20417 14047 20451
rect 16037 20417 16071 20451
rect 18981 20417 19015 20451
rect 21649 20417 21683 20451
rect 2145 20349 2179 20383
rect 6193 20349 6227 20383
rect 7205 20349 7239 20383
rect 7849 20349 7883 20383
rect 10701 20349 10735 20383
rect 13277 20349 13311 20383
rect 19625 20349 19659 20383
rect 9873 20281 9907 20315
rect 13645 20281 13679 20315
rect 14289 20281 14323 20315
rect 19349 20281 19383 20315
rect 19901 20281 19935 20315
rect 4537 20213 4571 20247
rect 4813 20213 4847 20247
rect 5825 20213 5859 20247
rect 11253 20213 11287 20247
rect 12725 20213 12759 20247
rect 2145 20009 2179 20043
rect 14105 20009 14139 20043
rect 16681 20009 16715 20043
rect 21281 20009 21315 20043
rect 1685 19941 1719 19975
rect 2421 19941 2455 19975
rect 5825 19941 5859 19975
rect 18981 19941 19015 19975
rect 22569 19941 22603 19975
rect 2513 19873 2547 19907
rect 4813 19873 4847 19907
rect 6101 19873 6135 19907
rect 9965 19873 9999 19907
rect 11529 19873 11563 19907
rect 12909 19873 12943 19907
rect 15577 19873 15611 19907
rect 17049 19873 17083 19907
rect 17233 19873 17267 19907
rect 17785 19873 17819 19907
rect 17969 19873 18003 19907
rect 19349 19873 19383 19907
rect 21097 19873 21131 19907
rect 22661 19873 22695 19907
rect 5273 19805 5307 19839
rect 6377 19805 6411 19839
rect 8125 19805 8159 19839
rect 11345 19805 11379 19839
rect 15485 19805 15519 19839
rect 16037 19805 16071 19839
rect 19257 19805 19291 19839
rect 3525 19669 3559 19703
rect 9321 19669 9355 19703
rect 10333 19669 10367 19703
rect 13093 19669 13127 19703
rect 14473 19669 14507 19703
rect 18245 19669 18279 19703
rect 21557 19669 21591 19703
rect 3801 19465 3835 19499
rect 4997 19465 5031 19499
rect 6285 19465 6319 19499
rect 8033 19465 8067 19499
rect 9137 19465 9171 19499
rect 16773 19465 16807 19499
rect 20913 19465 20947 19499
rect 22109 19465 22143 19499
rect 22753 19465 22787 19499
rect 9689 19397 9723 19431
rect 4445 19329 4479 19363
rect 5457 19329 5491 19363
rect 10701 19329 10735 19363
rect 17693 19329 17727 19363
rect 18521 19329 18555 19363
rect 20269 19329 20303 19363
rect 1685 19261 1719 19295
rect 2513 19261 2547 19295
rect 5365 19261 5399 19295
rect 5733 19261 5767 19295
rect 5917 19261 5951 19295
rect 7021 19261 7055 19295
rect 7665 19261 7699 19295
rect 8677 19261 8711 19295
rect 8953 19261 8987 19295
rect 10609 19261 10643 19295
rect 10977 19261 11011 19295
rect 11161 19261 11195 19295
rect 12081 19261 12115 19295
rect 12909 19261 12943 19295
rect 13737 19261 13771 19295
rect 15301 19261 15335 19295
rect 15577 19261 15611 19295
rect 16589 19261 16623 19295
rect 18245 19261 18279 19295
rect 21925 19261 21959 19295
rect 22385 19261 22419 19295
rect 11529 19193 11563 19227
rect 10057 19125 10091 19159
rect 15761 19125 15795 19159
rect 16037 19125 16071 19159
rect 17141 19125 17175 19159
rect 1685 18921 1719 18955
rect 4445 18921 4479 18955
rect 6561 18921 6595 18955
rect 7757 18921 7791 18955
rect 9321 18921 9355 18955
rect 10057 18921 10091 18955
rect 14473 18921 14507 18955
rect 16589 18921 16623 18955
rect 17509 18921 17543 18955
rect 18153 18921 18187 18955
rect 19257 18921 19291 18955
rect 19533 18921 19567 18955
rect 2421 18853 2455 18887
rect 7113 18853 7147 18887
rect 12725 18853 12759 18887
rect 17141 18853 17175 18887
rect 23121 18853 23155 18887
rect 1961 18785 1995 18819
rect 2973 18785 3007 18819
rect 5503 18785 5537 18819
rect 6101 18785 6135 18819
rect 6285 18785 6319 18819
rect 7573 18785 7607 18819
rect 15945 18785 15979 18819
rect 19073 18785 19107 18819
rect 5365 18717 5399 18751
rect 10701 18717 10735 18751
rect 10977 18717 11011 18751
rect 16221 18717 16255 18751
rect 19993 18717 20027 18751
rect 21097 18717 21131 18751
rect 21373 18717 21407 18751
rect 3157 18581 3191 18615
rect 4813 18581 4847 18615
rect 10333 18581 10367 18615
rect 13001 18581 13035 18615
rect 13461 18581 13495 18615
rect 18429 18581 18463 18615
rect 20545 18581 20579 18615
rect 5089 18377 5123 18411
rect 5733 18377 5767 18411
rect 7205 18377 7239 18411
rect 9229 18377 9263 18411
rect 21465 18377 21499 18411
rect 21741 18377 21775 18411
rect 5457 18309 5491 18343
rect 10977 18309 11011 18343
rect 11529 18309 11563 18343
rect 18429 18309 18463 18343
rect 2237 18241 2271 18275
rect 6101 18241 6135 18275
rect 7573 18241 7607 18275
rect 9597 18241 9631 18275
rect 14473 18241 14507 18275
rect 16497 18241 16531 18275
rect 16773 18241 16807 18275
rect 7021 18173 7055 18207
rect 7849 18173 7883 18207
rect 9873 18173 9907 18207
rect 10057 18173 10091 18207
rect 10517 18173 10551 18207
rect 10609 18173 10643 18207
rect 18245 18173 18279 18207
rect 18705 18173 18739 18207
rect 19625 18173 19659 18207
rect 20453 18173 20487 18207
rect 22293 18173 22327 18207
rect 22753 18173 22787 18207
rect 1961 18105 1995 18139
rect 2513 18105 2547 18139
rect 4261 18105 4295 18139
rect 4537 18105 4571 18139
rect 8861 18105 8895 18139
rect 14197 18105 14231 18139
rect 14749 18105 14783 18139
rect 8033 18037 8067 18071
rect 8309 18037 8343 18071
rect 19073 18037 19107 18071
rect 22477 18037 22511 18071
rect 2329 17833 2363 17867
rect 4445 17833 4479 17867
rect 8033 17833 8067 17867
rect 8677 17833 8711 17867
rect 9321 17833 9355 17867
rect 10793 17833 10827 17867
rect 14565 17833 14599 17867
rect 18981 17833 19015 17867
rect 19625 17833 19659 17867
rect 20453 17833 20487 17867
rect 2605 17765 2639 17799
rect 3065 17765 3099 17799
rect 13093 17765 13127 17799
rect 13921 17765 13955 17799
rect 14933 17765 14967 17799
rect 3341 17697 3375 17731
rect 4261 17697 4295 17731
rect 6377 17697 6411 17731
rect 7113 17697 7147 17731
rect 8493 17697 8527 17731
rect 9873 17697 9907 17731
rect 11529 17697 11563 17731
rect 12633 17697 12667 17731
rect 16129 17697 16163 17731
rect 16497 17697 16531 17731
rect 17693 17697 17727 17731
rect 18797 17697 18831 17731
rect 19257 17697 19291 17731
rect 4813 17629 4847 17663
rect 7481 17629 7515 17663
rect 12541 17629 12575 17663
rect 15485 17629 15519 17663
rect 15945 17629 15979 17663
rect 16405 17629 16439 17663
rect 18245 17629 18279 17663
rect 21465 17629 21499 17663
rect 21741 17629 21775 17663
rect 23489 17629 23523 17663
rect 1685 17493 1719 17527
rect 5365 17493 5399 17527
rect 10057 17493 10091 17527
rect 10333 17493 10367 17527
rect 11069 17493 11103 17527
rect 11713 17493 11747 17527
rect 17049 17493 17083 17527
rect 17417 17493 17451 17527
rect 17877 17493 17911 17527
rect 21097 17493 21131 17527
rect 6101 17289 6135 17323
rect 13277 17289 13311 17323
rect 15577 17289 15611 17323
rect 16497 17289 16531 17323
rect 17325 17289 17359 17323
rect 22569 17289 22603 17323
rect 13001 17221 13035 17255
rect 14933 17221 14967 17255
rect 20637 17221 20671 17255
rect 22017 17221 22051 17255
rect 1869 17153 1903 17187
rect 2421 17153 2455 17187
rect 17693 17153 17727 17187
rect 18521 17153 18555 17187
rect 20913 17153 20947 17187
rect 2145 17085 2179 17119
rect 4997 17085 5031 17119
rect 5365 17085 5399 17119
rect 6469 17085 6503 17119
rect 7113 17085 7147 17119
rect 9413 17085 9447 17119
rect 10057 17085 10091 17119
rect 12817 17085 12851 17119
rect 14013 17085 14047 17119
rect 14105 17085 14139 17119
rect 14473 17085 14507 17119
rect 14565 17085 14599 17119
rect 16681 17085 16715 17119
rect 18245 17085 18279 17119
rect 21097 17085 21131 17119
rect 21557 17085 21591 17119
rect 21649 17085 21683 17119
rect 4169 17017 4203 17051
rect 7021 17017 7055 17051
rect 20269 17017 20303 17051
rect 4537 16949 4571 16983
rect 8585 16949 8619 16983
rect 9045 16949 9079 16983
rect 11529 16949 11563 16983
rect 12081 16949 12115 16983
rect 22937 16949 22971 16983
rect 2237 16745 2271 16779
rect 3249 16745 3283 16779
rect 3709 16745 3743 16779
rect 6837 16745 6871 16779
rect 7297 16745 7331 16779
rect 9321 16745 9355 16779
rect 13553 16745 13587 16779
rect 14197 16745 14231 16779
rect 14841 16745 14875 16779
rect 17877 16745 17911 16779
rect 18613 16745 18647 16779
rect 19257 16745 19291 16779
rect 2881 16677 2915 16711
rect 4813 16677 4847 16711
rect 11069 16677 11103 16711
rect 13921 16677 13955 16711
rect 17509 16677 17543 16711
rect 20177 16677 20211 16711
rect 21649 16677 21683 16711
rect 5365 16609 5399 16643
rect 5457 16609 5491 16643
rect 5917 16609 5951 16643
rect 6101 16609 6135 16643
rect 8585 16609 8619 16643
rect 9873 16609 9907 16643
rect 15485 16609 15519 16643
rect 19073 16609 19107 16643
rect 22293 16609 22327 16643
rect 22661 16609 22695 16643
rect 1685 16541 1719 16575
rect 10793 16541 10827 16575
rect 12817 16541 12851 16575
rect 15761 16541 15795 16575
rect 22385 16541 22419 16575
rect 22569 16541 22603 16575
rect 6285 16473 6319 16507
rect 18337 16473 18371 16507
rect 2513 16405 2547 16439
rect 4353 16405 4387 16439
rect 8769 16405 8803 16439
rect 10057 16405 10091 16439
rect 13185 16405 13219 16439
rect 20545 16405 20579 16439
rect 21189 16405 21223 16439
rect 4997 16201 5031 16235
rect 6193 16201 6227 16235
rect 9873 16201 9907 16235
rect 10241 16201 10275 16235
rect 12817 16201 12851 16235
rect 15117 16201 15151 16235
rect 15853 16201 15887 16235
rect 16497 16201 16531 16235
rect 16589 16201 16623 16235
rect 16865 16201 16899 16235
rect 21005 16201 21039 16235
rect 22477 16201 22511 16235
rect 4077 16065 4111 16099
rect 7481 16065 7515 16099
rect 10517 16065 10551 16099
rect 15485 16065 15519 16099
rect 21373 16133 21407 16167
rect 21741 16065 21775 16099
rect 1685 15997 1719 16031
rect 2329 15997 2363 16031
rect 4445 15997 4479 16031
rect 5181 15997 5215 16031
rect 5365 15997 5399 16031
rect 5733 15997 5767 16031
rect 5825 15997 5859 16031
rect 7205 15997 7239 16031
rect 9229 15997 9263 16031
rect 10609 15997 10643 16031
rect 11069 15997 11103 16031
rect 12633 15997 12667 16031
rect 13093 15997 13127 16031
rect 14105 15997 14139 16031
rect 14565 15997 14599 16031
rect 16313 15997 16347 16031
rect 16589 15997 16623 16031
rect 18245 15997 18279 16031
rect 20637 15997 20671 16031
rect 22661 15997 22695 16031
rect 11345 15929 11379 15963
rect 18521 15929 18555 15963
rect 20269 15929 20303 15963
rect 11713 15861 11747 15895
rect 14289 15861 14323 15895
rect 17693 15861 17727 15895
rect 23121 15861 23155 15895
rect 7297 15657 7331 15691
rect 8585 15657 8619 15691
rect 10793 15657 10827 15691
rect 11161 15657 11195 15691
rect 18613 15657 18647 15691
rect 3249 15589 3283 15623
rect 4905 15589 4939 15623
rect 6653 15589 6687 15623
rect 16957 15589 16991 15623
rect 22569 15589 22603 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 2513 15521 2547 15555
rect 10241 15521 10275 15555
rect 13093 15521 13127 15555
rect 15945 15521 15979 15555
rect 18429 15521 18463 15555
rect 19533 15521 19567 15555
rect 21281 15521 21315 15555
rect 22661 15521 22695 15555
rect 1685 15453 1719 15487
rect 4629 15453 4663 15487
rect 7573 15453 7607 15487
rect 15853 15453 15887 15487
rect 19441 15453 19475 15487
rect 21189 15453 21223 15487
rect 2697 15385 2731 15419
rect 20269 15385 20303 15419
rect 22017 15385 22051 15419
rect 3617 15317 3651 15351
rect 4353 15317 4387 15351
rect 10425 15317 10459 15351
rect 12541 15317 12575 15351
rect 13185 15317 13219 15351
rect 14565 15317 14599 15351
rect 18153 15317 18187 15351
rect 19165 15317 19199 15351
rect 19717 15317 19751 15351
rect 21465 15317 21499 15351
rect 4721 15113 4755 15147
rect 6285 15113 6319 15147
rect 10241 15113 10275 15147
rect 15577 15113 15611 15147
rect 17693 15113 17727 15147
rect 20545 15113 20579 15147
rect 21925 15113 21959 15147
rect 22845 15113 22879 15147
rect 5273 15045 5307 15079
rect 11713 15045 11747 15079
rect 1961 14977 1995 15011
rect 2513 14977 2547 15011
rect 8493 14977 8527 15011
rect 9045 14977 9079 15011
rect 12081 14977 12115 15011
rect 13093 14977 13127 15011
rect 13553 14977 13587 15011
rect 14473 14977 14507 15011
rect 2237 14909 2271 14943
rect 5089 14909 5123 14943
rect 6009 14909 6043 14943
rect 7481 14909 7515 14943
rect 8585 14909 8619 14943
rect 9321 14909 9355 14943
rect 13277 14909 13311 14943
rect 13645 14909 13679 14943
rect 14197 14909 14231 14943
rect 14565 14909 14599 14943
rect 17049 14909 17083 14943
rect 18429 14909 18463 14943
rect 18889 14909 18923 14943
rect 20913 14909 20947 14943
rect 22385 14909 22419 14943
rect 23213 14909 23247 14943
rect 4261 14841 4295 14875
rect 7113 14841 7147 14875
rect 16405 14841 16439 14875
rect 20821 14841 20855 14875
rect 5549 14773 5583 14807
rect 7665 14773 7699 14807
rect 8033 14773 8067 14807
rect 12725 14773 12759 14807
rect 15945 14773 15979 14807
rect 22569 14773 22603 14807
rect 1869 14569 1903 14603
rect 3157 14569 3191 14603
rect 5641 14569 5675 14603
rect 8493 14569 8527 14603
rect 13185 14569 13219 14603
rect 13369 14569 13403 14603
rect 14381 14569 14415 14603
rect 19809 14569 19843 14603
rect 4077 14501 4111 14535
rect 4261 14501 4295 14535
rect 14933 14501 14967 14535
rect 23397 14501 23431 14535
rect 2237 14433 2271 14467
rect 2605 14433 2639 14467
rect 4905 14433 4939 14467
rect 7573 14433 7607 14467
rect 7941 14433 7975 14467
rect 10057 14433 10091 14467
rect 14197 14433 14231 14467
rect 15485 14433 15519 14467
rect 18797 14433 18831 14467
rect 19349 14433 19383 14467
rect 19533 14433 19567 14467
rect 2329 14365 2363 14399
rect 2513 14365 2547 14399
rect 3433 14365 3467 14399
rect 4077 14365 4111 14399
rect 7665 14365 7699 14399
rect 7849 14365 7883 14399
rect 11069 14365 11103 14399
rect 11345 14365 11379 14399
rect 15761 14365 15795 14399
rect 17509 14365 17543 14399
rect 18153 14365 18187 14399
rect 18613 14365 18647 14399
rect 21373 14365 21407 14399
rect 21649 14365 21683 14399
rect 6653 14297 6687 14331
rect 10701 14297 10735 14331
rect 6285 14229 6319 14263
rect 7205 14229 7239 14263
rect 10241 14229 10275 14263
rect 20453 14229 20487 14263
rect 1777 14025 1811 14059
rect 4997 14025 5031 14059
rect 9321 14025 9355 14059
rect 11437 14025 11471 14059
rect 14473 14025 14507 14059
rect 17693 14025 17727 14059
rect 20821 14025 20855 14059
rect 5733 13957 5767 13991
rect 6101 13957 6135 13991
rect 10701 13957 10735 13991
rect 11161 13957 11195 13991
rect 13737 13957 13771 13991
rect 22477 13957 22511 13991
rect 2697 13889 2731 13923
rect 7021 13889 7055 13923
rect 9045 13889 9079 13923
rect 9689 13889 9723 13923
rect 14841 13889 14875 13923
rect 15945 13889 15979 13923
rect 18797 13889 18831 13923
rect 19533 13889 19567 13923
rect 21097 13889 21131 13923
rect 22845 13889 22879 13923
rect 1593 13821 1627 13855
rect 5549 13821 5583 13855
rect 9781 13821 9815 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 13369 13821 13403 13855
rect 13553 13821 13587 13855
rect 16129 13821 16163 13855
rect 16497 13821 16531 13855
rect 16589 13821 16623 13855
rect 18429 13821 18463 13855
rect 19717 13821 19751 13855
rect 20085 13821 20119 13855
rect 20269 13821 20303 13855
rect 21649 13821 21683 13855
rect 2421 13753 2455 13787
rect 2973 13753 3007 13787
rect 4721 13753 4755 13787
rect 6469 13753 6503 13787
rect 7297 13753 7331 13787
rect 12081 13753 12115 13787
rect 17325 13753 17359 13787
rect 19073 13753 19107 13787
rect 15209 13685 15243 13719
rect 15577 13685 15611 13719
rect 22109 13685 22143 13719
rect 2605 13481 2639 13515
rect 8309 13481 8343 13515
rect 9229 13481 9263 13515
rect 12541 13481 12575 13515
rect 14197 13481 14231 13515
rect 16681 13481 16715 13515
rect 17141 13481 17175 13515
rect 19165 13481 19199 13515
rect 19441 13481 19475 13515
rect 19809 13481 19843 13515
rect 3249 13413 3283 13447
rect 6837 13413 6871 13447
rect 10149 13413 10183 13447
rect 11897 13413 11931 13447
rect 13185 13413 13219 13447
rect 14933 13413 14967 13447
rect 17785 13413 17819 13447
rect 20545 13413 20579 13447
rect 2789 13345 2823 13379
rect 4629 13345 4663 13379
rect 5181 13345 5215 13379
rect 7113 13345 7147 13379
rect 7297 13345 7331 13379
rect 7849 13345 7883 13379
rect 8033 13345 8067 13379
rect 15669 13345 15703 13379
rect 16129 13345 16163 13379
rect 16221 13345 16255 13379
rect 18429 13345 18463 13379
rect 21557 13345 21591 13379
rect 21741 13345 21775 13379
rect 9873 13277 9907 13311
rect 15485 13277 15519 13311
rect 1593 13141 1627 13175
rect 3525 13141 3559 13175
rect 12817 13141 12851 13175
rect 18153 13141 18187 13175
rect 18613 13141 18647 13175
rect 2421 12937 2455 12971
rect 3157 12937 3191 12971
rect 4445 12937 4479 12971
rect 4813 12937 4847 12971
rect 5549 12937 5583 12971
rect 8309 12937 8343 12971
rect 10149 12937 10183 12971
rect 16405 12937 16439 12971
rect 16773 12937 16807 12971
rect 17233 12937 17267 12971
rect 3433 12869 3467 12903
rect 8677 12869 8711 12903
rect 2145 12801 2179 12835
rect 1593 12733 1627 12767
rect 1685 12733 1719 12767
rect 2881 12665 2915 12699
rect 6469 12801 6503 12835
rect 7297 12801 7331 12835
rect 20269 12801 20303 12835
rect 5365 12733 5399 12767
rect 5825 12733 5859 12767
rect 7389 12733 7423 12767
rect 13921 12733 13955 12767
rect 14381 12733 14415 12767
rect 15117 12733 15151 12767
rect 18245 12733 18279 12767
rect 20729 12733 20763 12767
rect 21005 12733 21039 12767
rect 21741 12733 21775 12767
rect 22109 12733 22143 12767
rect 9321 12665 9355 12699
rect 11161 12665 11195 12699
rect 11989 12665 12023 12699
rect 12725 12665 12759 12699
rect 13093 12665 13127 12699
rect 17693 12665 17727 12699
rect 18521 12665 18555 12699
rect 22017 12665 22051 12699
rect 3433 12597 3467 12631
rect 3525 12597 3559 12631
rect 9781 12597 9815 12631
rect 10517 12597 10551 12631
rect 11253 12597 11287 12631
rect 21189 12597 21223 12631
rect 2513 12393 2547 12427
rect 2789 12393 2823 12427
rect 5365 12393 5399 12427
rect 7389 12393 7423 12427
rect 7757 12393 7791 12427
rect 8217 12393 8251 12427
rect 12633 12393 12667 12427
rect 14473 12393 14507 12427
rect 15485 12393 15519 12427
rect 16313 12393 16347 12427
rect 17693 12393 17727 12427
rect 19993 12393 20027 12427
rect 20545 12325 20579 12359
rect 23397 12325 23431 12359
rect 1685 12257 1719 12291
rect 4905 12257 4939 12291
rect 8033 12257 8067 12291
rect 10149 12257 10183 12291
rect 10517 12257 10551 12291
rect 11345 12257 11379 12291
rect 13185 12257 13219 12291
rect 14013 12257 14047 12291
rect 15853 12257 15887 12291
rect 18429 12257 18463 12291
rect 18797 12257 18831 12291
rect 19257 12257 19291 12291
rect 19809 12257 19843 12291
rect 21373 12257 21407 12291
rect 1593 12189 1627 12223
rect 2145 12189 2179 12223
rect 13645 12189 13679 12223
rect 21649 12189 21683 12223
rect 13369 12121 13403 12155
rect 18153 12121 18187 12155
rect 3157 12053 3191 12087
rect 3617 12053 3651 12087
rect 5089 12053 5123 12087
rect 14933 12053 14967 12087
rect 16037 12053 16071 12087
rect 18981 12053 19015 12087
rect 1685 11849 1719 11883
rect 7021 11849 7055 11883
rect 10517 11849 10551 11883
rect 12817 11849 12851 11883
rect 13921 11849 13955 11883
rect 9229 11781 9263 11815
rect 9505 11781 9539 11815
rect 21097 11781 21131 11815
rect 22477 11781 22511 11815
rect 3617 11713 3651 11747
rect 5641 11713 5675 11747
rect 7941 11713 7975 11747
rect 10241 11713 10275 11747
rect 13645 11713 13679 11747
rect 15025 11713 15059 11747
rect 15301 11713 15335 11747
rect 18245 11713 18279 11747
rect 2697 11645 2731 11679
rect 8585 11645 8619 11679
rect 9505 11645 9539 11679
rect 9597 11645 9631 11679
rect 9689 11645 9723 11679
rect 10977 11645 11011 11679
rect 11069 11645 11103 11679
rect 12633 11645 12667 11679
rect 13093 11645 13127 11679
rect 13737 11645 13771 11679
rect 21557 11645 21591 11679
rect 21649 11645 21683 11679
rect 22017 11645 22051 11679
rect 22109 11645 22143 11679
rect 3341 11577 3375 11611
rect 3893 11577 3927 11611
rect 8309 11577 8343 11611
rect 10149 11577 10183 11611
rect 10241 11577 10275 11611
rect 11529 11577 11563 11611
rect 17049 11577 17083 11611
rect 17693 11577 17727 11611
rect 18521 11577 18555 11611
rect 20269 11577 20303 11611
rect 23029 11577 23063 11611
rect 2513 11509 2547 11543
rect 8769 11509 8803 11543
rect 11897 11509 11931 11543
rect 14565 11509 14599 11543
rect 20637 11509 20671 11543
rect 23857 11509 23891 11543
rect 2421 11305 2455 11339
rect 10057 11305 10091 11339
rect 10425 11305 10459 11339
rect 14933 11305 14967 11339
rect 21281 11305 21315 11339
rect 21649 11305 21683 11339
rect 3709 11237 3743 11271
rect 12541 11237 12575 11271
rect 13461 11237 13495 11271
rect 15945 11237 15979 11271
rect 16865 11237 16899 11271
rect 20545 11237 20579 11271
rect 1593 11169 1627 11203
rect 5641 11169 5675 11203
rect 6101 11169 6135 11203
rect 7573 11169 7607 11203
rect 9873 11169 9907 11203
rect 10793 11169 10827 11203
rect 14565 11169 14599 11203
rect 15485 11169 15519 11203
rect 17417 11169 17451 11203
rect 18061 11169 18095 11203
rect 21097 11169 21131 11203
rect 22017 11169 22051 11203
rect 22477 11169 22511 11203
rect 22661 11169 22695 11203
rect 23029 11169 23063 11203
rect 7021 11101 7055 11135
rect 22937 11101 22971 11135
rect 1777 11033 1811 11067
rect 13645 11033 13679 11067
rect 15669 11033 15703 11067
rect 20177 11033 20211 11067
rect 2053 10965 2087 10999
rect 2881 10965 2915 10999
rect 3249 10965 3283 10999
rect 4261 10965 4295 10999
rect 7757 10965 7791 10999
rect 6009 10761 6043 10795
rect 10793 10761 10827 10795
rect 11897 10761 11931 10795
rect 13461 10761 13495 10795
rect 14105 10761 14139 10795
rect 14749 10761 14783 10795
rect 22017 10761 22051 10795
rect 22385 10761 22419 10795
rect 23029 10761 23063 10795
rect 19349 10693 19383 10727
rect 5089 10625 5123 10659
rect 7021 10625 7055 10659
rect 9413 10625 9447 10659
rect 14473 10625 14507 10659
rect 22661 10625 22695 10659
rect 1869 10557 1903 10591
rect 2513 10557 2547 10591
rect 3893 10557 3927 10591
rect 4629 10557 4663 10591
rect 4813 10557 4847 10591
rect 5181 10557 5215 10591
rect 9689 10557 9723 10591
rect 11161 10557 11195 10591
rect 12633 10557 12667 10591
rect 13093 10557 13127 10591
rect 14565 10557 14599 10591
rect 16129 10557 16163 10591
rect 16865 10557 16899 10591
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 18981 10557 19015 10591
rect 19165 10557 19199 10591
rect 20269 10557 20303 10591
rect 20361 10557 20395 10591
rect 21833 10557 21867 10591
rect 3525 10489 3559 10523
rect 4169 10489 4203 10523
rect 6469 10489 6503 10523
rect 7297 10489 7331 10523
rect 9045 10489 9079 10523
rect 17141 10489 17175 10523
rect 23857 10489 23891 10523
rect 5641 10421 5675 10455
rect 9873 10421 9907 10455
rect 10241 10421 10275 10455
rect 11253 10421 11287 10455
rect 12817 10421 12851 10455
rect 15393 10421 15427 10455
rect 15761 10421 15795 10455
rect 17693 10421 17727 10455
rect 19901 10421 19935 10455
rect 21281 10421 21315 10455
rect 3525 10217 3559 10251
rect 5641 10217 5675 10251
rect 7297 10217 7331 10251
rect 8493 10217 8527 10251
rect 10425 10217 10459 10251
rect 13829 10217 13863 10251
rect 17601 10217 17635 10251
rect 21281 10217 21315 10251
rect 21557 10217 21591 10251
rect 22017 10217 22051 10251
rect 23029 10217 23063 10251
rect 5365 10149 5399 10183
rect 17049 10149 17083 10183
rect 1961 10081 1995 10115
rect 2513 10081 2547 10115
rect 2697 10081 2731 10115
rect 4261 10081 4295 10115
rect 4721 10081 4755 10115
rect 6285 10081 6319 10115
rect 6377 10081 6411 10115
rect 6837 10081 6871 10115
rect 7021 10081 7055 10115
rect 8309 10081 8343 10115
rect 10241 10081 10275 10115
rect 12909 10081 12943 10115
rect 13093 10081 13127 10115
rect 15577 10081 15611 10115
rect 16681 10081 16715 10115
rect 17969 10081 18003 10115
rect 18337 10081 18371 10115
rect 18797 10081 18831 10115
rect 21097 10081 21131 10115
rect 22661 10081 22695 10115
rect 1869 10013 1903 10047
rect 12173 10013 12207 10047
rect 15485 10013 15519 10047
rect 17785 10013 17819 10047
rect 18245 10013 18279 10047
rect 8769 9945 8803 9979
rect 12541 9945 12575 9979
rect 2973 9877 3007 9911
rect 7757 9877 7791 9911
rect 9965 9877 9999 9911
rect 13185 9877 13219 9911
rect 14933 9877 14967 9911
rect 15761 9877 15795 9911
rect 2053 9673 2087 9707
rect 5365 9673 5399 9707
rect 8493 9673 8527 9707
rect 16865 9673 16899 9707
rect 17417 9673 17451 9707
rect 18613 9673 18647 9707
rect 20361 9673 20395 9707
rect 22477 9673 22511 9707
rect 23857 9673 23891 9707
rect 6101 9605 6135 9639
rect 18337 9605 18371 9639
rect 2421 9537 2455 9571
rect 2973 9537 3007 9571
rect 4721 9537 4755 9571
rect 7021 9537 7055 9571
rect 7941 9537 7975 9571
rect 12081 9537 12115 9571
rect 12909 9537 12943 9571
rect 2697 9469 2731 9503
rect 6469 9469 6503 9503
rect 7481 9469 7515 9503
rect 7665 9469 7699 9503
rect 8033 9469 8067 9503
rect 10149 9469 10183 9503
rect 10885 9469 10919 9503
rect 11253 9469 11287 9503
rect 12633 9469 12667 9503
rect 14933 9469 14967 9503
rect 15301 9469 15335 9503
rect 15393 9469 15427 9503
rect 16681 9469 16715 9503
rect 20177 9469 20211 9503
rect 20637 9469 20671 9503
rect 22201 9469 22235 9503
rect 22293 9469 22327 9503
rect 9505 9401 9539 9435
rect 11621 9401 11655 9435
rect 14657 9401 14691 9435
rect 15853 9401 15887 9435
rect 19073 9401 19107 9435
rect 1685 9333 1719 9367
rect 5733 9333 5767 9367
rect 9229 9333 9263 9367
rect 10609 9333 10643 9367
rect 16129 9333 16163 9367
rect 21097 9333 21131 9367
rect 21833 9333 21867 9367
rect 23121 9333 23155 9367
rect 3433 9129 3467 9163
rect 4261 9129 4295 9163
rect 5825 9129 5859 9163
rect 6193 9129 6227 9163
rect 9321 9129 9355 9163
rect 9965 9129 9999 9163
rect 14933 9129 14967 9163
rect 17785 9129 17819 9163
rect 3157 9061 3191 9095
rect 6929 9061 6963 9095
rect 17417 9061 17451 9095
rect 23489 9061 23523 9095
rect 1685 8993 1719 9027
rect 5089 8993 5123 9027
rect 7021 8993 7055 9027
rect 8585 8993 8619 9027
rect 10517 8993 10551 9027
rect 10885 8993 10919 9027
rect 11345 8993 11379 9027
rect 12265 8993 12299 9027
rect 13001 8993 13035 9027
rect 15577 8993 15611 9027
rect 18613 8993 18647 9027
rect 1593 8925 1627 8959
rect 10333 8925 10367 8959
rect 10793 8925 10827 8959
rect 13277 8925 13311 8959
rect 15485 8925 15519 8959
rect 16681 8925 16715 8959
rect 21465 8925 21499 8959
rect 21741 8925 21775 8959
rect 2789 8857 2823 8891
rect 4721 8857 4755 8891
rect 6653 8857 6687 8891
rect 12541 8857 12575 8891
rect 18245 8857 18279 8891
rect 1869 8789 1903 8823
rect 5273 8789 5307 8823
rect 7941 8789 7975 8823
rect 8769 8789 8803 8823
rect 15761 8789 15795 8823
rect 18797 8789 18831 8823
rect 19533 8789 19567 8823
rect 2053 8585 2087 8619
rect 3525 8585 3559 8619
rect 4058 8585 4092 8619
rect 9413 8585 9447 8619
rect 12817 8585 12851 8619
rect 13093 8585 13127 8619
rect 16405 8585 16439 8619
rect 20821 8585 20855 8619
rect 21833 8585 21867 8619
rect 3157 8449 3191 8483
rect 7021 8449 7055 8483
rect 9045 8449 9079 8483
rect 15485 8449 15519 8483
rect 20269 8449 20303 8483
rect 21557 8449 21591 8483
rect 1593 8381 1627 8415
rect 3801 8381 3835 8415
rect 5825 8381 5859 8415
rect 9689 8381 9723 8415
rect 9873 8381 9907 8415
rect 10425 8381 10459 8415
rect 10609 8381 10643 8415
rect 12633 8381 12667 8415
rect 14381 8381 14415 8415
rect 15853 8381 15887 8415
rect 16681 8381 16715 8415
rect 18245 8381 18279 8415
rect 21649 8381 21683 8415
rect 6469 8313 6503 8347
rect 7297 8313 7331 8347
rect 17233 8313 17267 8347
rect 17693 8313 17727 8347
rect 18521 8313 18555 8347
rect 22477 8313 22511 8347
rect 1777 8245 1811 8279
rect 2513 8245 2547 8279
rect 10885 8245 10919 8279
rect 11345 8245 11379 8279
rect 11989 8245 12023 8279
rect 14013 8245 14047 8279
rect 14749 8245 14783 8279
rect 16037 8245 16071 8279
rect 21281 8245 21315 8279
rect 22753 8245 22787 8279
rect 3433 8041 3467 8075
rect 4445 8041 4479 8075
rect 5089 8041 5123 8075
rect 5917 8041 5951 8075
rect 7297 8041 7331 8075
rect 7941 8041 7975 8075
rect 9321 8041 9355 8075
rect 12357 8041 12391 8075
rect 12725 8041 12759 8075
rect 21281 8041 21315 8075
rect 21649 8041 21683 8075
rect 22293 8041 22327 8075
rect 22569 8041 22603 8075
rect 8309 7973 8343 8007
rect 10149 7973 10183 8007
rect 16221 7973 16255 8007
rect 2421 7905 2455 7939
rect 4261 7905 4295 7939
rect 6837 7905 6871 7939
rect 7757 7905 7791 7939
rect 8585 7905 8619 7939
rect 14933 7905 14967 7939
rect 15485 7905 15519 7939
rect 16589 7905 16623 7939
rect 17417 7905 17451 7939
rect 19349 7905 19383 7939
rect 21097 7905 21131 7939
rect 22109 7905 22143 7939
rect 23121 7905 23155 7939
rect 9873 7837 9907 7871
rect 11897 7837 11931 7871
rect 18429 7837 18463 7871
rect 19257 7837 19291 7871
rect 20269 7769 20303 7803
rect 1593 7701 1627 7735
rect 2053 7701 2087 7735
rect 2605 7701 2639 7735
rect 6653 7701 6687 7735
rect 14105 7701 14139 7735
rect 15669 7701 15703 7735
rect 18705 7701 18739 7735
rect 23305 7701 23339 7735
rect 7481 7497 7515 7531
rect 10149 7497 10183 7531
rect 20453 7497 20487 7531
rect 23213 7497 23247 7531
rect 7205 7429 7239 7463
rect 19349 7429 19383 7463
rect 2881 7361 2915 7395
rect 11345 7361 11379 7395
rect 14105 7361 14139 7395
rect 16313 7361 16347 7395
rect 18245 7361 18279 7395
rect 1685 7293 1719 7327
rect 2421 7293 2455 7327
rect 2605 7293 2639 7327
rect 2973 7293 3007 7327
rect 4077 7293 4111 7327
rect 6285 7293 6319 7327
rect 8769 7293 8803 7327
rect 9229 7293 9263 7327
rect 10701 7293 10735 7327
rect 14289 7293 14323 7327
rect 14749 7293 14783 7327
rect 14841 7293 14875 7327
rect 16405 7293 16439 7327
rect 18429 7293 18463 7327
rect 18889 7293 18923 7327
rect 18981 7293 19015 7327
rect 20085 7293 20119 7327
rect 20821 7293 20855 7327
rect 21557 7293 21591 7327
rect 1961 7225 1995 7259
rect 13829 7225 13863 7259
rect 17693 7225 17727 7259
rect 3525 7157 3559 7191
rect 4261 7157 4295 7191
rect 4629 7157 4663 7191
rect 4997 7157 5031 7191
rect 13369 7157 13403 7191
rect 15301 7157 15335 7191
rect 15945 7157 15979 7191
rect 3617 6953 3651 6987
rect 9965 6953 9999 6987
rect 14197 6953 14231 6987
rect 14841 6953 14875 6987
rect 16957 6953 16991 6987
rect 17969 6953 18003 6987
rect 4537 6885 4571 6919
rect 10241 6885 10275 6919
rect 10609 6885 10643 6919
rect 11897 6885 11931 6919
rect 15485 6885 15519 6919
rect 17417 6885 17451 6919
rect 20545 6885 20579 6919
rect 1777 6817 1811 6851
rect 2237 6817 2271 6851
rect 2329 6817 2363 6851
rect 5457 6817 5491 6851
rect 6193 6817 6227 6851
rect 7941 6817 7975 6851
rect 11621 6817 11655 6851
rect 13645 6817 13679 6851
rect 14565 6817 14599 6851
rect 16129 6817 16163 6851
rect 16497 6817 16531 6851
rect 18337 6817 18371 6851
rect 18659 6817 18693 6851
rect 18797 6817 18831 6851
rect 19809 6817 19843 6851
rect 1685 6749 1719 6783
rect 15945 6749 15979 6783
rect 16405 6749 16439 6783
rect 18153 6749 18187 6783
rect 21557 6749 21591 6783
rect 21833 6749 21867 6783
rect 23581 6749 23615 6783
rect 2697 6681 2731 6715
rect 3249 6613 3283 6647
rect 7113 6613 7147 6647
rect 7849 6613 7883 6647
rect 19165 6613 19199 6647
rect 19993 6613 20027 6647
rect 21281 6613 21315 6647
rect 1777 6409 1811 6443
rect 4905 6409 4939 6443
rect 11897 6409 11931 6443
rect 12633 6409 12667 6443
rect 17325 6409 17359 6443
rect 17693 6409 17727 6443
rect 21097 6409 21131 6443
rect 22569 6409 22603 6443
rect 23121 6409 23155 6443
rect 5825 6341 5859 6375
rect 11069 6341 11103 6375
rect 11529 6341 11563 6375
rect 2145 6273 2179 6307
rect 2697 6273 2731 6307
rect 4445 6273 4479 6307
rect 7941 6273 7975 6307
rect 14473 6273 14507 6307
rect 15025 6273 15059 6307
rect 16773 6273 16807 6307
rect 18429 6273 18463 6307
rect 18705 6273 18739 6307
rect 21373 6273 21407 6307
rect 2421 6205 2455 6239
rect 5273 6205 5307 6239
rect 7481 6205 7515 6239
rect 7665 6205 7699 6239
rect 8033 6205 8067 6239
rect 8861 6205 8895 6239
rect 9965 6205 9999 6239
rect 10425 6205 10459 6239
rect 11345 6205 11379 6239
rect 14105 6205 14139 6239
rect 14749 6205 14783 6239
rect 21557 6205 21591 6239
rect 22109 6205 22143 6239
rect 22293 6205 22327 6239
rect 7021 6137 7055 6171
rect 20453 6137 20487 6171
rect 23857 6137 23891 6171
rect 5457 6069 5491 6103
rect 6469 6069 6503 6103
rect 8585 6069 8619 6103
rect 9045 6069 9079 6103
rect 9413 6069 9447 6103
rect 10149 6069 10183 6103
rect 1685 5865 1719 5899
rect 3433 5865 3467 5899
rect 6653 5865 6687 5899
rect 8585 5865 8619 5899
rect 10149 5865 10183 5899
rect 11805 5865 11839 5899
rect 15577 5865 15611 5899
rect 15945 5865 15979 5899
rect 16681 5865 16715 5899
rect 17785 5865 17819 5899
rect 18521 5865 18555 5899
rect 19257 5865 19291 5899
rect 20545 5865 20579 5899
rect 21925 5865 21959 5899
rect 23121 5865 23155 5899
rect 2053 5797 2087 5831
rect 3157 5797 3191 5831
rect 6285 5797 6319 5831
rect 17049 5797 17083 5831
rect 17417 5797 17451 5831
rect 19901 5797 19935 5831
rect 2605 5729 2639 5763
rect 7113 5729 7147 5763
rect 7573 5729 7607 5763
rect 7665 5729 7699 5763
rect 9965 5729 9999 5763
rect 11345 5729 11379 5763
rect 13001 5729 13035 5763
rect 13737 5729 13771 5763
rect 19073 5729 19107 5763
rect 22293 5729 22327 5763
rect 22661 5729 22695 5763
rect 22845 5729 22879 5763
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 6929 5661 6963 5695
rect 22385 5661 22419 5695
rect 8033 5593 8067 5627
rect 11529 5593 11563 5627
rect 18153 5593 18187 5627
rect 14749 5525 14783 5559
rect 21373 5525 21407 5559
rect 4537 5321 4571 5355
rect 5365 5321 5399 5355
rect 6469 5321 6503 5355
rect 11069 5321 11103 5355
rect 11713 5321 11747 5355
rect 12725 5321 12759 5355
rect 21465 5321 21499 5355
rect 22017 5321 22051 5355
rect 4169 5253 4203 5287
rect 4813 5253 4847 5287
rect 6101 5253 6135 5287
rect 13921 5253 13955 5287
rect 21097 5253 21131 5287
rect 5733 5185 5767 5219
rect 7205 5185 7239 5219
rect 7757 5185 7791 5219
rect 9505 5185 9539 5219
rect 17693 5185 17727 5219
rect 18521 5185 18555 5219
rect 20269 5185 20303 5219
rect 1685 5117 1719 5151
rect 2237 5117 2271 5151
rect 7481 5117 7515 5151
rect 10885 5117 10919 5151
rect 13093 5117 13127 5151
rect 13553 5117 13587 5151
rect 15117 5117 15151 5151
rect 16221 5117 16255 5151
rect 16681 5117 16715 5151
rect 17141 5117 17175 5151
rect 18245 5117 18279 5151
rect 21833 5117 21867 5151
rect 22753 5117 22787 5151
rect 14473 5049 14507 5083
rect 15577 5049 15611 5083
rect 10057 4981 10091 5015
rect 11345 4981 11379 5015
rect 13277 4981 13311 5015
rect 15853 4981 15887 5015
rect 16865 4981 16899 5015
rect 1685 4777 1719 4811
rect 2053 4777 2087 4811
rect 2329 4777 2363 4811
rect 3065 4777 3099 4811
rect 3433 4777 3467 4811
rect 4813 4777 4847 4811
rect 7849 4777 7883 4811
rect 12357 4777 12391 4811
rect 18429 4777 18463 4811
rect 21373 4777 21407 4811
rect 22017 4777 22051 4811
rect 8125 4709 8159 4743
rect 13553 4709 13587 4743
rect 18797 4709 18831 4743
rect 21741 4709 21775 4743
rect 22845 4709 22879 4743
rect 4261 4641 4295 4675
rect 5917 4641 5951 4675
rect 6009 4641 6043 4675
rect 6377 4641 6411 4675
rect 6469 4641 6503 4675
rect 8585 4641 8619 4675
rect 9873 4641 9907 4675
rect 11345 4641 11379 4675
rect 13001 4641 13035 4675
rect 18245 4641 18279 4675
rect 19073 4641 19107 4675
rect 21189 4641 21223 4675
rect 23489 4641 23523 4675
rect 7021 4573 7055 4607
rect 7389 4573 7423 4607
rect 14565 4573 14599 4607
rect 15485 4573 15519 4607
rect 15761 4573 15795 4607
rect 17509 4573 17543 4607
rect 22385 4573 22419 4607
rect 10057 4505 10091 4539
rect 11529 4505 11563 4539
rect 14841 4505 14875 4539
rect 4445 4437 4479 4471
rect 5365 4437 5399 4471
rect 8769 4437 8803 4471
rect 12725 4437 12759 4471
rect 13185 4437 13219 4471
rect 17969 4437 18003 4471
rect 20177 4437 20211 4471
rect 20545 4437 20579 4471
rect 2605 4233 2639 4267
rect 5457 4233 5491 4267
rect 9781 4233 9815 4267
rect 10885 4233 10919 4267
rect 17141 4233 17175 4267
rect 17601 4233 17635 4267
rect 22477 4233 22511 4267
rect 22937 4233 22971 4267
rect 15209 4165 15243 4199
rect 16589 4165 16623 4199
rect 3249 4097 3283 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 12633 4097 12667 4131
rect 12909 4097 12943 4131
rect 14657 4097 14691 4131
rect 21925 4097 21959 4131
rect 2973 4029 3007 4063
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 16129 4029 16163 4063
rect 16221 4029 16255 4063
rect 19165 4029 19199 4063
rect 19625 4029 19659 4063
rect 20729 4029 20763 4063
rect 21465 4029 21499 4063
rect 21649 4029 21683 4063
rect 22017 4029 22051 4063
rect 4997 3961 5031 3995
rect 6469 3961 6503 3995
rect 9229 3961 9263 3995
rect 11529 3961 11563 3995
rect 5733 3893 5767 3927
rect 10241 3893 10275 3927
rect 11805 3893 11839 3927
rect 21281 3893 21315 3927
rect 3065 3689 3099 3723
rect 4813 3689 4847 3723
rect 12725 3689 12759 3723
rect 14933 3689 14967 3723
rect 19993 3689 20027 3723
rect 8493 3621 8527 3655
rect 10517 3621 10551 3655
rect 12265 3621 12299 3655
rect 16221 3621 16255 3655
rect 3709 3553 3743 3587
rect 5181 3553 5215 3587
rect 5549 3553 5583 3587
rect 5733 3553 5767 3587
rect 6653 3553 6687 3587
rect 7205 3553 7239 3587
rect 13829 3553 13863 3587
rect 14197 3553 14231 3587
rect 14381 3553 14415 3587
rect 16037 3553 16071 3587
rect 16957 3553 16991 3587
rect 19809 3553 19843 3587
rect 20269 3553 20303 3587
rect 4997 3485 5031 3519
rect 10241 3485 10275 3519
rect 13645 3485 13679 3519
rect 17233 3485 17267 3519
rect 18981 3485 19015 3519
rect 21097 3485 21131 3519
rect 21373 3485 21407 3519
rect 23121 3485 23155 3519
rect 6009 3349 6043 3383
rect 8861 3349 8895 3383
rect 13461 3349 13495 3383
rect 19533 3349 19567 3383
rect 9873 3145 9907 3179
rect 10885 3145 10919 3179
rect 11437 3145 11471 3179
rect 12909 3145 12943 3179
rect 13553 3145 13587 3179
rect 16129 3145 16163 3179
rect 16681 3145 16715 3179
rect 17417 3145 17451 3179
rect 21925 3145 21959 3179
rect 22661 3145 22695 3179
rect 8125 3077 8159 3111
rect 21373 3077 21407 3111
rect 22293 3077 22327 3111
rect 2053 3009 2087 3043
rect 4629 3009 4663 3043
rect 7021 3009 7055 3043
rect 9321 3009 9355 3043
rect 9597 3009 9631 3043
rect 15761 3009 15795 3043
rect 16957 3009 16991 3043
rect 19441 3009 19475 3043
rect 20361 3009 20395 3043
rect 2145 2941 2179 2975
rect 3525 2941 3559 2975
rect 4169 2941 4203 2975
rect 5457 2941 5491 2975
rect 7665 2941 7699 2975
rect 9689 2941 9723 2975
rect 11253 2941 11287 2975
rect 11989 2941 12023 2975
rect 12633 2941 12667 2975
rect 12725 2941 12759 2975
rect 14749 2941 14783 2975
rect 15209 2941 15243 2975
rect 18889 2941 18923 2975
rect 18981 2941 19015 2975
rect 20453 2941 20487 2975
rect 20919 2941 20953 2975
rect 21005 2941 21039 2975
rect 2605 2873 2639 2907
rect 5181 2873 5215 2907
rect 10517 2873 10551 2907
rect 19809 2873 19843 2907
rect 23029 2873 23063 2907
rect 1685 2805 1719 2839
rect 3065 2805 3099 2839
rect 6377 2805 6411 2839
rect 18521 2805 18555 2839
rect 2053 2601 2087 2635
rect 3617 2601 3651 2635
rect 4169 2601 4203 2635
rect 4445 2601 4479 2635
rect 4813 2601 4847 2635
rect 5457 2601 5491 2635
rect 7113 2601 7147 2635
rect 7573 2601 7607 2635
rect 10241 2601 10275 2635
rect 10609 2601 10643 2635
rect 11253 2601 11287 2635
rect 11897 2601 11931 2635
rect 13277 2601 13311 2635
rect 13737 2601 13771 2635
rect 14105 2601 14139 2635
rect 14473 2601 14507 2635
rect 18705 2601 18739 2635
rect 19073 2601 19107 2635
rect 19993 2601 20027 2635
rect 20637 2601 20671 2635
rect 21373 2601 21407 2635
rect 21741 2601 21775 2635
rect 5089 2533 5123 2567
rect 14749 2533 14783 2567
rect 22109 2533 22143 2567
rect 12265 2465 12299 2499
rect 12817 2465 12851 2499
rect 18521 2465 18555 2499
rect 19625 2465 19659 2499
rect 22201 2465 22235 2499
rect 17969 2397 18003 2431
rect 13001 2329 13035 2363
<< metal1 >>
rect 8386 27208 8392 27260
rect 8444 27248 8450 27260
rect 11698 27248 11704 27260
rect 8444 27220 11704 27248
rect 8444 27208 8450 27220
rect 11698 27208 11704 27220
rect 11756 27208 11762 27260
rect 1104 25594 24656 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 24656 25594
rect 1104 25520 24656 25542
rect 4982 25344 4988 25356
rect 4895 25316 4988 25344
rect 4982 25304 4988 25316
rect 5040 25344 5046 25356
rect 5534 25344 5540 25356
rect 5040 25316 5540 25344
rect 5040 25304 5046 25316
rect 5534 25304 5540 25316
rect 5592 25304 5598 25356
rect 8386 25344 8392 25356
rect 8347 25316 8392 25344
rect 8386 25304 8392 25316
rect 8444 25304 8450 25356
rect 12253 25347 12311 25353
rect 12253 25313 12265 25347
rect 12299 25344 12311 25347
rect 12618 25344 12624 25356
rect 12299 25316 12624 25344
rect 12299 25313 12311 25316
rect 12253 25307 12311 25313
rect 12618 25304 12624 25316
rect 12676 25344 12682 25356
rect 13081 25347 13139 25353
rect 13081 25344 13093 25347
rect 12676 25316 13093 25344
rect 12676 25304 12682 25316
rect 13081 25313 13093 25316
rect 13127 25313 13139 25347
rect 13081 25307 13139 25313
rect 13170 25304 13176 25356
rect 13228 25344 13234 25356
rect 15657 25347 15715 25353
rect 15657 25344 15669 25347
rect 13228 25316 15669 25344
rect 13228 25304 13234 25316
rect 15657 25313 15669 25316
rect 15703 25344 15715 25347
rect 16114 25344 16120 25356
rect 15703 25316 16120 25344
rect 15703 25313 15715 25316
rect 15657 25307 15715 25313
rect 16114 25304 16120 25316
rect 16172 25304 16178 25356
rect 16758 25344 16764 25356
rect 16719 25316 16764 25344
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 22373 25347 22431 25353
rect 22373 25313 22385 25347
rect 22419 25344 22431 25347
rect 22462 25344 22468 25356
rect 22419 25316 22468 25344
rect 22419 25313 22431 25316
rect 22373 25307 22431 25313
rect 22462 25304 22468 25316
rect 22520 25344 22526 25356
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22520 25316 22845 25344
rect 22520 25304 22526 25316
rect 22833 25313 22845 25316
rect 22879 25313 22891 25347
rect 22833 25307 22891 25313
rect 2038 25236 2044 25288
rect 2096 25276 2102 25288
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 2096 25248 4905 25276
rect 2096 25236 2102 25248
rect 4893 25245 4905 25248
rect 4939 25276 4951 25279
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 4939 25248 5733 25276
rect 4939 25245 4951 25248
rect 4893 25239 4951 25245
rect 5721 25245 5733 25248
rect 5767 25276 5779 25279
rect 7282 25276 7288 25288
rect 5767 25248 7288 25276
rect 5767 25245 5779 25248
rect 5721 25239 5779 25245
rect 7282 25236 7288 25248
rect 7340 25276 7346 25288
rect 8297 25279 8355 25285
rect 8297 25276 8309 25279
rect 7340 25248 8309 25276
rect 7340 25236 7346 25248
rect 8297 25245 8309 25248
rect 8343 25245 8355 25279
rect 8297 25239 8355 25245
rect 14093 25211 14151 25217
rect 14093 25177 14105 25211
rect 14139 25208 14151 25211
rect 14182 25208 14188 25220
rect 14139 25180 14188 25208
rect 14139 25177 14151 25180
rect 14093 25171 14151 25177
rect 14182 25168 14188 25180
rect 14240 25208 14246 25220
rect 15841 25211 15899 25217
rect 15841 25208 15853 25211
rect 14240 25180 15853 25208
rect 14240 25168 14246 25180
rect 15841 25177 15853 25180
rect 15887 25177 15899 25211
rect 15841 25171 15899 25177
rect 5166 25140 5172 25152
rect 5127 25112 5172 25140
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 8570 25140 8576 25152
rect 8531 25112 8576 25140
rect 8570 25100 8576 25112
rect 8628 25100 8634 25152
rect 9398 25100 9404 25152
rect 9456 25140 9462 25152
rect 10045 25143 10103 25149
rect 10045 25140 10057 25143
rect 9456 25112 10057 25140
rect 9456 25100 9462 25112
rect 10045 25109 10057 25112
rect 10091 25140 10103 25143
rect 10410 25140 10416 25152
rect 10091 25112 10416 25140
rect 10091 25109 10103 25112
rect 10045 25103 10103 25109
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 10870 25140 10876 25152
rect 10831 25112 10876 25140
rect 10870 25100 10876 25112
rect 10928 25100 10934 25152
rect 13449 25143 13507 25149
rect 13449 25109 13461 25143
rect 13495 25140 13507 25143
rect 13538 25140 13544 25152
rect 13495 25112 13544 25140
rect 13495 25109 13507 25112
rect 13449 25103 13507 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 14458 25140 14464 25152
rect 14419 25112 14464 25140
rect 14458 25100 14464 25112
rect 14516 25100 14522 25152
rect 16942 25140 16948 25152
rect 16903 25112 16948 25140
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 22554 25140 22560 25152
rect 22515 25112 22560 25140
rect 22554 25100 22560 25112
rect 22612 25100 22618 25152
rect 1104 25050 24656 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 24656 25050
rect 1104 24976 24656 24998
rect 4893 24939 4951 24945
rect 4893 24905 4905 24939
rect 4939 24936 4951 24939
rect 4982 24936 4988 24948
rect 4939 24908 4988 24936
rect 4939 24905 4951 24908
rect 4893 24899 4951 24905
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 7282 24936 7288 24948
rect 7243 24908 7288 24936
rect 7282 24896 7288 24908
rect 7340 24896 7346 24948
rect 8294 24936 8300 24948
rect 8255 24908 8300 24936
rect 8294 24896 8300 24908
rect 8352 24896 8358 24948
rect 16114 24936 16120 24948
rect 9646 24908 10548 24936
rect 16075 24908 16120 24936
rect 9646 24868 9674 24908
rect 8128 24840 9674 24868
rect 10520 24868 10548 24908
rect 16114 24896 16120 24908
rect 16172 24896 16178 24948
rect 16758 24936 16764 24948
rect 16719 24908 16764 24936
rect 16758 24896 16764 24908
rect 16816 24896 16822 24948
rect 22462 24936 22468 24948
rect 22423 24908 22468 24936
rect 22462 24896 22468 24908
rect 22520 24896 22526 24948
rect 23106 24936 23112 24948
rect 23067 24908 23112 24936
rect 23106 24896 23112 24908
rect 23164 24896 23170 24948
rect 25498 24868 25504 24880
rect 10520 24840 25504 24868
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24800 7803 24803
rect 8128 24800 8156 24840
rect 25498 24828 25504 24840
rect 25556 24828 25562 24880
rect 9398 24800 9404 24812
rect 7791 24772 8156 24800
rect 9359 24772 9404 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24732 3939 24735
rect 4157 24735 4215 24741
rect 4157 24732 4169 24735
rect 3927 24704 4169 24732
rect 3927 24701 3939 24704
rect 3881 24695 3939 24701
rect 4157 24701 4169 24704
rect 4203 24732 4215 24735
rect 5166 24732 5172 24744
rect 4203 24704 5172 24732
rect 4203 24701 4215 24704
rect 4157 24695 4215 24701
rect 5166 24692 5172 24704
rect 5224 24692 5230 24744
rect 5813 24735 5871 24741
rect 5813 24701 5825 24735
rect 5859 24732 5871 24735
rect 6181 24735 6239 24741
rect 6181 24732 6193 24735
rect 5859 24704 6193 24732
rect 5859 24701 5871 24704
rect 5813 24695 5871 24701
rect 6181 24701 6193 24704
rect 6227 24732 6239 24735
rect 6362 24732 6368 24744
rect 6227 24704 6368 24732
rect 6227 24701 6239 24704
rect 6181 24695 6239 24701
rect 6362 24692 6368 24704
rect 6420 24692 6426 24744
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7558 24732 7564 24744
rect 7340 24704 7564 24732
rect 7340 24692 7346 24704
rect 7558 24692 7564 24704
rect 7616 24732 7622 24744
rect 8018 24732 8024 24744
rect 7616 24704 8024 24732
rect 7616 24692 7622 24704
rect 8018 24692 8024 24704
rect 8076 24692 8082 24744
rect 8128 24741 8156 24772
rect 9398 24760 9404 24772
rect 9456 24760 9462 24812
rect 10410 24760 10416 24812
rect 10468 24800 10474 24812
rect 11054 24800 11060 24812
rect 10468 24772 11060 24800
rect 10468 24760 10474 24772
rect 11054 24760 11060 24772
rect 11112 24800 11118 24812
rect 12621 24803 12679 24809
rect 12621 24800 12633 24803
rect 11112 24772 12633 24800
rect 11112 24760 11118 24772
rect 12621 24769 12633 24772
rect 12667 24800 12679 24803
rect 13170 24800 13176 24812
rect 12667 24772 12940 24800
rect 13131 24772 13176 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 8113 24735 8171 24741
rect 8113 24701 8125 24735
rect 8159 24701 8171 24735
rect 8113 24695 8171 24701
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24732 9551 24735
rect 10321 24735 10379 24741
rect 10321 24732 10333 24735
rect 9539 24704 10333 24732
rect 9539 24701 9551 24704
rect 9493 24695 9551 24701
rect 10321 24701 10333 24704
rect 10367 24732 10379 24735
rect 10594 24732 10600 24744
rect 10367 24704 10600 24732
rect 10367 24701 10379 24704
rect 10321 24695 10379 24701
rect 10594 24692 10600 24704
rect 10652 24692 10658 24744
rect 10870 24732 10876 24744
rect 10831 24704 10876 24732
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 12713 24735 12771 24741
rect 12713 24701 12725 24735
rect 12759 24701 12771 24735
rect 12912 24732 12940 24772
rect 13170 24760 13176 24772
rect 13228 24760 13234 24812
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 12912 24704 13461 24732
rect 12713 24695 12771 24701
rect 13449 24701 13461 24704
rect 13495 24701 13507 24735
rect 14182 24732 14188 24744
rect 14143 24704 14188 24732
rect 13449 24695 13507 24701
rect 9858 24624 9864 24676
rect 9916 24664 9922 24676
rect 9953 24667 10011 24673
rect 9953 24664 9965 24667
rect 9916 24636 9965 24664
rect 9916 24624 9922 24636
rect 9953 24633 9965 24636
rect 9999 24633 10011 24667
rect 11514 24664 11520 24676
rect 11475 24636 11520 24664
rect 9953 24627 10011 24633
rect 11514 24624 11520 24636
rect 11572 24624 11578 24676
rect 12069 24667 12127 24673
rect 12069 24633 12081 24667
rect 12115 24664 12127 24667
rect 12728 24664 12756 24695
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14458 24692 14464 24744
rect 14516 24732 14522 24744
rect 14553 24735 14611 24741
rect 14553 24732 14565 24735
rect 14516 24704 14565 24732
rect 14516 24692 14522 24704
rect 14553 24701 14565 24704
rect 14599 24701 14611 24735
rect 15930 24732 15936 24744
rect 14553 24695 14611 24701
rect 14844 24704 15936 24732
rect 14844 24664 14872 24704
rect 15930 24692 15936 24704
rect 15988 24692 15994 24744
rect 18874 24732 18880 24744
rect 18835 24704 18880 24732
rect 18874 24692 18880 24704
rect 18932 24692 18938 24744
rect 18966 24692 18972 24744
rect 19024 24732 19030 24744
rect 19613 24735 19671 24741
rect 19613 24732 19625 24735
rect 19024 24704 19625 24732
rect 19024 24692 19030 24704
rect 19613 24701 19625 24704
rect 19659 24732 19671 24735
rect 20901 24735 20959 24741
rect 19659 24704 19932 24732
rect 19659 24701 19671 24704
rect 19613 24695 19671 24701
rect 12115 24636 14872 24664
rect 12115 24633 12127 24636
rect 12069 24627 12127 24633
rect 14918 24624 14924 24676
rect 14976 24624 14982 24676
rect 17681 24667 17739 24673
rect 17681 24633 17693 24667
rect 17727 24664 17739 24667
rect 18984 24664 19012 24692
rect 17727 24636 19012 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 4341 24599 4399 24605
rect 4341 24565 4353 24599
rect 4387 24596 4399 24599
rect 4706 24596 4712 24608
rect 4387 24568 4712 24596
rect 4387 24565 4399 24568
rect 4341 24559 4399 24565
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5350 24556 5356 24608
rect 5408 24596 5414 24608
rect 5445 24599 5503 24605
rect 5445 24596 5457 24599
rect 5408 24568 5457 24596
rect 5408 24556 5414 24568
rect 5445 24565 5457 24568
rect 5491 24565 5503 24599
rect 5445 24559 5503 24565
rect 8386 24556 8392 24608
rect 8444 24596 8450 24608
rect 8941 24599 8999 24605
rect 8941 24596 8953 24599
rect 8444 24568 8953 24596
rect 8444 24556 8450 24568
rect 8941 24565 8953 24568
rect 8987 24596 8999 24599
rect 13078 24596 13084 24608
rect 8987 24568 13084 24596
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 13078 24556 13084 24568
rect 13136 24556 13142 24608
rect 17310 24596 17316 24608
rect 17271 24568 17316 24596
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 18690 24556 18696 24608
rect 18748 24596 18754 24608
rect 19260 24596 19288 24664
rect 18748 24568 19288 24596
rect 19904 24596 19932 24704
rect 20901 24701 20913 24735
rect 20947 24732 20959 24735
rect 21177 24735 21235 24741
rect 21177 24732 21189 24735
rect 20947 24704 21189 24732
rect 20947 24701 20959 24704
rect 20901 24695 20959 24701
rect 21177 24701 21189 24704
rect 21223 24732 21235 24735
rect 21450 24732 21456 24744
rect 21223 24704 21456 24732
rect 21223 24701 21235 24704
rect 21177 24695 21235 24701
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 22189 24735 22247 24741
rect 22189 24732 22201 24735
rect 21836 24704 22201 24732
rect 21361 24599 21419 24605
rect 21361 24596 21373 24599
rect 19904 24568 21373 24596
rect 18748 24556 18754 24568
rect 21361 24565 21373 24568
rect 21407 24565 21419 24599
rect 21361 24559 21419 24565
rect 21726 24556 21732 24608
rect 21784 24596 21790 24608
rect 21836 24605 21864 24704
rect 22189 24701 22201 24704
rect 22235 24701 22247 24735
rect 22189 24695 22247 24701
rect 22281 24735 22339 24741
rect 22281 24701 22293 24735
rect 22327 24732 22339 24735
rect 23106 24732 23112 24744
rect 22327 24704 23112 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 23106 24692 23112 24704
rect 23164 24692 23170 24744
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21784 24568 21833 24596
rect 21784 24556 21790 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 1104 24506 24656 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 24656 24506
rect 1104 24432 24656 24454
rect 8018 24352 8024 24404
rect 8076 24392 8082 24404
rect 9033 24395 9091 24401
rect 9033 24392 9045 24395
rect 8076 24364 9045 24392
rect 8076 24352 8082 24364
rect 9033 24361 9045 24364
rect 9079 24361 9091 24395
rect 9033 24355 9091 24361
rect 14182 24352 14188 24404
rect 14240 24392 14246 24404
rect 14829 24395 14887 24401
rect 14829 24392 14841 24395
rect 14240 24364 14841 24392
rect 14240 24352 14246 24364
rect 14829 24361 14841 24364
rect 14875 24392 14887 24395
rect 15470 24392 15476 24404
rect 14875 24364 15476 24392
rect 14875 24361 14887 24364
rect 14829 24355 14887 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 17310 24352 17316 24404
rect 17368 24392 17374 24404
rect 17865 24395 17923 24401
rect 17865 24392 17877 24395
rect 17368 24364 17877 24392
rect 17368 24352 17374 24364
rect 17865 24361 17877 24364
rect 17911 24392 17923 24395
rect 18874 24392 18880 24404
rect 17911 24364 18880 24392
rect 17911 24361 17923 24364
rect 17865 24355 17923 24361
rect 3326 24284 3332 24336
rect 3384 24324 3390 24336
rect 3384 24296 8340 24324
rect 3384 24284 3390 24296
rect 1670 24256 1676 24268
rect 1631 24228 1676 24256
rect 1670 24216 1676 24228
rect 1728 24216 1734 24268
rect 4614 24256 4620 24268
rect 4575 24228 4620 24256
rect 4614 24216 4620 24228
rect 4672 24216 4678 24268
rect 4706 24216 4712 24268
rect 4764 24256 4770 24268
rect 5166 24256 5172 24268
rect 4764 24228 4809 24256
rect 5127 24228 5172 24256
rect 4764 24216 4770 24228
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 5350 24256 5356 24268
rect 5311 24228 5356 24256
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 6365 24259 6423 24265
rect 6365 24225 6377 24259
rect 6411 24256 6423 24259
rect 6733 24259 6791 24265
rect 6733 24256 6745 24259
rect 6411 24228 6745 24256
rect 6411 24225 6423 24228
rect 6365 24219 6423 24225
rect 6733 24225 6745 24228
rect 6779 24256 6791 24259
rect 7650 24256 7656 24268
rect 6779 24228 7656 24256
rect 6779 24225 6791 24228
rect 6733 24219 6791 24225
rect 7650 24216 7656 24228
rect 7708 24216 7714 24268
rect 8312 24265 8340 24296
rect 14458 24284 14464 24336
rect 14516 24324 14522 24336
rect 15654 24324 15660 24336
rect 14516 24296 15660 24324
rect 14516 24284 14522 24296
rect 15654 24284 15660 24296
rect 15712 24324 15718 24336
rect 15749 24327 15807 24333
rect 15749 24324 15761 24327
rect 15712 24296 15761 24324
rect 15712 24284 15718 24296
rect 15749 24293 15761 24296
rect 15795 24324 15807 24327
rect 17221 24327 17279 24333
rect 17221 24324 17233 24327
rect 15795 24296 17233 24324
rect 15795 24293 15807 24296
rect 15749 24287 15807 24293
rect 17221 24293 17233 24296
rect 17267 24293 17279 24327
rect 17221 24287 17279 24293
rect 8297 24259 8355 24265
rect 8297 24225 8309 24259
rect 8343 24256 8355 24259
rect 8478 24256 8484 24268
rect 8343 24228 8484 24256
rect 8343 24225 8355 24228
rect 8297 24219 8355 24225
rect 8478 24216 8484 24228
rect 8536 24216 8542 24268
rect 10962 24256 10968 24268
rect 10923 24228 10968 24256
rect 10962 24216 10968 24228
rect 11020 24216 11026 24268
rect 11422 24256 11428 24268
rect 11335 24228 11428 24256
rect 11422 24216 11428 24228
rect 11480 24256 11486 24268
rect 11480 24228 11652 24256
rect 11480 24216 11486 24228
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 2038 24188 2044 24200
rect 1627 24160 2044 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 2958 24148 2964 24200
rect 3016 24188 3022 24200
rect 4724 24188 4752 24216
rect 3016 24160 4752 24188
rect 7377 24191 7435 24197
rect 3016 24148 3022 24160
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 7742 24188 7748 24200
rect 7423 24160 7748 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7742 24148 7748 24160
rect 7800 24148 7806 24200
rect 8205 24191 8263 24197
rect 8205 24157 8217 24191
rect 8251 24157 8263 24191
rect 8754 24188 8760 24200
rect 8715 24160 8760 24188
rect 8205 24151 8263 24157
rect 4982 24080 4988 24132
rect 5040 24120 5046 24132
rect 5537 24123 5595 24129
rect 5537 24120 5549 24123
rect 5040 24092 5549 24120
rect 5040 24080 5046 24092
rect 5537 24089 5549 24092
rect 5583 24089 5595 24123
rect 8220 24120 8248 24151
rect 8754 24148 8760 24160
rect 8812 24148 8818 24200
rect 11624 24188 11652 24228
rect 12250 24216 12256 24268
rect 12308 24256 12314 24268
rect 12943 24259 13001 24265
rect 12943 24256 12955 24259
rect 12308 24228 12955 24256
rect 12308 24216 12314 24228
rect 12943 24225 12955 24228
rect 12989 24225 13001 24259
rect 13446 24256 13452 24268
rect 13407 24228 13452 24256
rect 12943 24219 13001 24225
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 14553 24259 14611 24265
rect 13596 24228 13641 24256
rect 13596 24216 13602 24228
rect 14553 24225 14565 24259
rect 14599 24256 14611 24259
rect 16298 24256 16304 24268
rect 14599 24228 16304 24256
rect 14599 24225 14611 24228
rect 14553 24219 14611 24225
rect 16298 24216 16304 24228
rect 16356 24256 16362 24268
rect 16393 24259 16451 24265
rect 16393 24256 16405 24259
rect 16356 24228 16405 24256
rect 16356 24216 16362 24228
rect 16393 24225 16405 24228
rect 16439 24225 16451 24259
rect 16758 24256 16764 24268
rect 16719 24228 16764 24256
rect 16393 24219 16451 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 16942 24256 16948 24268
rect 16903 24228 16948 24256
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 18800 24265 18828 24364
rect 18874 24352 18880 24364
rect 18932 24352 18938 24404
rect 22646 24352 22652 24404
rect 22704 24352 22710 24404
rect 19150 24284 19156 24336
rect 19208 24324 19214 24336
rect 19208 24296 19564 24324
rect 19208 24284 19214 24296
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24225 18843 24259
rect 18785 24219 18843 24225
rect 18877 24259 18935 24265
rect 18877 24225 18889 24259
rect 18923 24256 18935 24259
rect 18966 24256 18972 24268
rect 18923 24228 18972 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 12802 24188 12808 24200
rect 11624 24160 12808 24188
rect 12802 24148 12808 24160
rect 12860 24148 12866 24200
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 16666 24188 16672 24200
rect 16531 24160 16672 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 18325 24191 18383 24197
rect 18325 24157 18337 24191
rect 18371 24188 18383 24191
rect 18892 24188 18920 24219
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 19334 24216 19340 24268
rect 19392 24256 19398 24268
rect 19536 24265 19564 24296
rect 19521 24259 19579 24265
rect 19392 24228 19437 24256
rect 19392 24216 19398 24228
rect 19521 24225 19533 24259
rect 19567 24256 19579 24259
rect 21174 24256 21180 24268
rect 19567 24228 20392 24256
rect 21135 24228 21180 24256
rect 19567 24225 19579 24228
rect 19521 24219 19579 24225
rect 20364 24200 20392 24228
rect 21174 24216 21180 24228
rect 21232 24216 21238 24268
rect 22664 24265 22692 24352
rect 22649 24259 22707 24265
rect 22649 24225 22661 24259
rect 22695 24225 22707 24259
rect 22649 24219 22707 24225
rect 18371 24160 18920 24188
rect 18371 24157 18383 24160
rect 18325 24151 18383 24157
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 20404 24160 21097 24188
rect 20404 24148 20410 24160
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22557 24191 22615 24197
rect 22557 24188 22569 24191
rect 21784 24160 22569 24188
rect 21784 24148 21790 24160
rect 22557 24157 22569 24160
rect 22603 24188 22615 24191
rect 22922 24188 22928 24200
rect 22603 24160 22928 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 22922 24148 22928 24160
rect 22980 24148 22986 24200
rect 9398 24120 9404 24132
rect 8220 24092 9404 24120
rect 5537 24083 5595 24089
rect 9398 24080 9404 24092
rect 9456 24080 9462 24132
rect 12894 24080 12900 24132
rect 12952 24120 12958 24132
rect 13909 24123 13967 24129
rect 13909 24120 13921 24123
rect 12952 24092 13921 24120
rect 12952 24080 12958 24092
rect 13909 24089 13921 24092
rect 13955 24089 13967 24123
rect 13909 24083 13967 24089
rect 18506 24080 18512 24132
rect 18564 24120 18570 24132
rect 19705 24123 19763 24129
rect 19705 24120 19717 24123
rect 18564 24092 19717 24120
rect 18564 24080 18570 24092
rect 19705 24089 19717 24092
rect 19751 24089 19763 24123
rect 19705 24083 19763 24089
rect 1854 24052 1860 24064
rect 1815 24024 1860 24052
rect 1854 24012 1860 24024
rect 1912 24012 1918 24064
rect 2593 24055 2651 24061
rect 2593 24021 2605 24055
rect 2639 24052 2651 24055
rect 3142 24052 3148 24064
rect 2639 24024 3148 24052
rect 2639 24021 2651 24024
rect 2593 24015 2651 24021
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 11974 24052 11980 24064
rect 11935 24024 11980 24052
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 12342 24012 12348 24064
rect 12400 24052 12406 24064
rect 12437 24055 12495 24061
rect 12437 24052 12449 24055
rect 12400 24024 12449 24052
rect 12400 24012 12406 24024
rect 12437 24021 12449 24024
rect 12483 24021 12495 24055
rect 12437 24015 12495 24021
rect 21450 24012 21456 24064
rect 21508 24052 21514 24064
rect 22833 24055 22891 24061
rect 22833 24052 22845 24055
rect 21508 24024 22845 24052
rect 21508 24012 21514 24024
rect 22833 24021 22845 24024
rect 22879 24021 22891 24055
rect 22833 24015 22891 24021
rect 1104 23962 24656 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 24656 23962
rect 1104 23888 24656 23910
rect 1670 23848 1676 23860
rect 1631 23820 1676 23848
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 2038 23848 2044 23860
rect 1999 23820 2044 23848
rect 2038 23808 2044 23820
rect 2096 23808 2102 23860
rect 4801 23851 4859 23857
rect 4801 23817 4813 23851
rect 4847 23848 4859 23851
rect 5350 23848 5356 23860
rect 4847 23820 5356 23848
rect 4847 23817 4859 23820
rect 4801 23811 4859 23817
rect 5350 23808 5356 23820
rect 5408 23848 5414 23860
rect 5902 23848 5908 23860
rect 5408 23820 5908 23848
rect 5408 23808 5414 23820
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 6362 23848 6368 23860
rect 6323 23820 6368 23848
rect 6362 23808 6368 23820
rect 6420 23808 6426 23860
rect 8478 23848 8484 23860
rect 8439 23820 8484 23848
rect 8478 23808 8484 23820
rect 8536 23808 8542 23860
rect 8941 23851 8999 23857
rect 8941 23817 8953 23851
rect 8987 23848 8999 23851
rect 9398 23848 9404 23860
rect 8987 23820 9404 23848
rect 8987 23817 8999 23820
rect 8941 23811 8999 23817
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 9769 23851 9827 23857
rect 9769 23817 9781 23851
rect 9815 23848 9827 23851
rect 10505 23851 10563 23857
rect 10505 23848 10517 23851
rect 9815 23820 10517 23848
rect 9815 23817 9827 23820
rect 9769 23811 9827 23817
rect 10505 23817 10517 23820
rect 10551 23848 10563 23851
rect 11422 23848 11428 23860
rect 10551 23820 11428 23848
rect 10551 23817 10563 23820
rect 10505 23811 10563 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 11606 23808 11612 23860
rect 11664 23848 11670 23860
rect 11701 23851 11759 23857
rect 11701 23848 11713 23851
rect 11664 23820 11713 23848
rect 11664 23808 11670 23820
rect 11701 23817 11713 23820
rect 11747 23848 11759 23851
rect 13538 23848 13544 23860
rect 11747 23820 13544 23848
rect 11747 23817 11759 23820
rect 11701 23811 11759 23817
rect 13538 23808 13544 23820
rect 13596 23808 13602 23860
rect 15197 23851 15255 23857
rect 15197 23817 15209 23851
rect 15243 23848 15255 23851
rect 16666 23848 16672 23860
rect 15243 23820 16672 23848
rect 15243 23817 15255 23820
rect 15197 23811 15255 23817
rect 16666 23808 16672 23820
rect 16724 23808 16730 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17497 23851 17555 23857
rect 17497 23848 17509 23851
rect 16816 23820 17509 23848
rect 16816 23808 16822 23820
rect 17497 23817 17509 23820
rect 17543 23817 17555 23851
rect 17497 23811 17555 23817
rect 18877 23851 18935 23857
rect 18877 23817 18889 23851
rect 18923 23848 18935 23851
rect 20438 23848 20444 23860
rect 18923 23820 20444 23848
rect 18923 23817 18935 23820
rect 18877 23811 18935 23817
rect 4706 23740 4712 23792
rect 4764 23780 4770 23792
rect 5445 23783 5503 23789
rect 5445 23780 5457 23783
rect 4764 23752 5457 23780
rect 4764 23740 4770 23752
rect 5445 23749 5457 23752
rect 5491 23749 5503 23783
rect 5445 23743 5503 23749
rect 10873 23783 10931 23789
rect 10873 23749 10885 23783
rect 10919 23780 10931 23783
rect 10962 23780 10968 23792
rect 10919 23752 10968 23780
rect 10919 23749 10931 23752
rect 10873 23743 10931 23749
rect 10962 23740 10968 23752
rect 11020 23780 11026 23792
rect 11333 23783 11391 23789
rect 11333 23780 11345 23783
rect 11020 23752 11345 23780
rect 11020 23740 11026 23752
rect 11333 23749 11345 23752
rect 11379 23780 11391 23783
rect 12250 23780 12256 23792
rect 11379 23752 12256 23780
rect 11379 23749 11391 23752
rect 11333 23743 11391 23749
rect 12250 23740 12256 23752
rect 12308 23740 12314 23792
rect 16114 23740 16120 23792
rect 16172 23780 16178 23792
rect 16390 23780 16396 23792
rect 16172 23752 16396 23780
rect 16172 23740 16178 23752
rect 16390 23740 16396 23752
rect 16448 23780 16454 23792
rect 16942 23780 16948 23792
rect 16448 23752 16948 23780
rect 16448 23740 16454 23752
rect 16942 23740 16948 23752
rect 17000 23780 17006 23792
rect 17129 23783 17187 23789
rect 17129 23780 17141 23783
rect 17000 23752 17141 23780
rect 17000 23740 17006 23752
rect 17129 23749 17141 23752
rect 17175 23749 17187 23783
rect 17129 23743 17187 23749
rect 5166 23712 5172 23724
rect 5079 23684 5172 23712
rect 5166 23672 5172 23684
rect 5224 23712 5230 23724
rect 6089 23715 6147 23721
rect 6089 23712 6101 23715
rect 5224 23684 6101 23712
rect 5224 23672 5230 23684
rect 6089 23681 6101 23684
rect 6135 23712 6147 23715
rect 12069 23715 12127 23721
rect 6135 23684 7788 23712
rect 6135 23681 6147 23684
rect 6089 23675 6147 23681
rect 7760 23656 7788 23684
rect 12069 23681 12081 23715
rect 12115 23712 12127 23715
rect 12894 23712 12900 23724
rect 12115 23684 12900 23712
rect 12115 23681 12127 23684
rect 12069 23675 12127 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 15470 23712 15476 23724
rect 15431 23684 15476 23712
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 18874 23672 18880 23724
rect 18932 23712 18938 23724
rect 19720 23721 19748 23820
rect 20438 23808 20444 23820
rect 20496 23848 20502 23860
rect 20901 23851 20959 23857
rect 20901 23848 20913 23851
rect 20496 23820 20913 23848
rect 20496 23808 20502 23820
rect 20901 23817 20913 23820
rect 20947 23848 20959 23851
rect 21174 23848 21180 23860
rect 20947 23820 21180 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 22646 23848 22652 23860
rect 22607 23820 22652 23848
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 22922 23848 22928 23860
rect 22883 23820 22928 23848
rect 22922 23808 22928 23820
rect 22980 23808 22986 23860
rect 19153 23715 19211 23721
rect 19153 23712 19165 23715
rect 18932 23684 19165 23712
rect 18932 23672 18938 23684
rect 19153 23681 19165 23684
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19978 23712 19984 23724
rect 19705 23675 19763 23681
rect 19812 23684 19984 23712
rect 2590 23604 2596 23656
rect 2648 23644 2654 23656
rect 2958 23644 2964 23656
rect 2648 23616 2964 23644
rect 2648 23604 2654 23616
rect 2958 23604 2964 23616
rect 3016 23604 3022 23656
rect 3142 23644 3148 23656
rect 3103 23616 3148 23644
rect 3142 23604 3148 23616
rect 3200 23644 3206 23656
rect 3200 23616 4660 23644
rect 3200 23604 3206 23616
rect 4632 23588 4660 23616
rect 6362 23604 6368 23656
rect 6420 23644 6426 23656
rect 7469 23647 7527 23653
rect 7469 23644 7481 23647
rect 6420 23616 7481 23644
rect 6420 23604 6426 23616
rect 7469 23613 7481 23616
rect 7515 23613 7527 23647
rect 7650 23644 7656 23656
rect 7611 23616 7656 23644
rect 7469 23607 7527 23613
rect 7650 23604 7656 23616
rect 7708 23604 7714 23656
rect 7742 23604 7748 23656
rect 7800 23644 7806 23656
rect 7975 23647 8033 23653
rect 7975 23644 7987 23647
rect 7800 23616 7987 23644
rect 7800 23604 7806 23616
rect 7975 23613 7987 23616
rect 8021 23613 8033 23647
rect 8110 23644 8116 23656
rect 8071 23616 8116 23644
rect 7975 23607 8033 23613
rect 8110 23604 8116 23616
rect 8168 23604 8174 23656
rect 8754 23604 8760 23656
rect 8812 23644 8818 23656
rect 9585 23647 9643 23653
rect 9585 23644 9597 23647
rect 8812 23616 9597 23644
rect 8812 23604 8818 23616
rect 9585 23613 9597 23616
rect 9631 23644 9643 23647
rect 10045 23647 10103 23653
rect 10045 23644 10057 23647
rect 9631 23616 10057 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 10045 23613 10057 23616
rect 10091 23613 10103 23647
rect 10045 23607 10103 23613
rect 12526 23604 12532 23656
rect 12584 23644 12590 23656
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12584 23616 12633 23644
rect 12584 23604 12590 23616
rect 12621 23613 12633 23616
rect 12667 23613 12679 23647
rect 15654 23644 15660 23656
rect 15615 23616 15660 23644
rect 12621 23607 12679 23613
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 16114 23644 16120 23656
rect 16075 23616 16120 23644
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 16209 23647 16267 23653
rect 16209 23613 16221 23647
rect 16255 23644 16267 23647
rect 16758 23644 16764 23656
rect 16255 23616 16764 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 2406 23536 2412 23588
rect 2464 23576 2470 23588
rect 2464 23548 3556 23576
rect 2464 23536 2470 23548
rect 4614 23536 4620 23588
rect 4672 23576 4678 23588
rect 7009 23579 7067 23585
rect 7009 23576 7021 23579
rect 4672 23548 7021 23576
rect 4672 23536 4678 23548
rect 7009 23545 7021 23548
rect 7055 23545 7067 23579
rect 7009 23539 7067 23545
rect 12342 23536 12348 23588
rect 12400 23576 12406 23588
rect 14642 23576 14648 23588
rect 12400 23548 13400 23576
rect 14603 23548 14648 23576
rect 12400 23536 12406 23548
rect 14642 23536 14648 23548
rect 14700 23536 14706 23588
rect 16022 23536 16028 23588
rect 16080 23576 16086 23588
rect 16224 23576 16252 23607
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 19812 23653 19840 23684
rect 19978 23672 19984 23684
rect 20036 23712 20042 23724
rect 20036 23684 21864 23712
rect 20036 23672 20042 23684
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 20162 23604 20168 23656
rect 20220 23644 20226 23656
rect 20346 23644 20352 23656
rect 20220 23616 20265 23644
rect 20307 23616 20352 23644
rect 20220 23604 20226 23616
rect 20346 23604 20352 23616
rect 20404 23604 20410 23656
rect 21836 23653 21864 23684
rect 21821 23647 21879 23653
rect 21821 23613 21833 23647
rect 21867 23644 21879 23647
rect 22189 23647 22247 23653
rect 22189 23644 22201 23647
rect 21867 23616 22201 23644
rect 21867 23613 21879 23616
rect 21821 23607 21879 23613
rect 22189 23613 22201 23616
rect 22235 23613 22247 23647
rect 22189 23607 22247 23613
rect 16080 23548 16252 23576
rect 18509 23579 18567 23585
rect 16080 23536 16086 23548
rect 18509 23545 18521 23579
rect 18555 23576 18567 23579
rect 19150 23576 19156 23588
rect 18555 23548 19156 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 19150 23536 19156 23548
rect 19208 23536 19214 23588
rect 21174 23576 21180 23588
rect 21135 23548 21180 23576
rect 21174 23536 21180 23548
rect 21232 23536 21238 23588
rect 16206 23468 16212 23520
rect 16264 23508 16270 23520
rect 16669 23511 16727 23517
rect 16669 23508 16681 23511
rect 16264 23480 16681 23508
rect 16264 23468 16270 23480
rect 16669 23477 16681 23480
rect 16715 23477 16727 23511
rect 16669 23471 16727 23477
rect 1104 23418 24656 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 24656 23418
rect 1104 23344 24656 23366
rect 2590 23304 2596 23316
rect 2551 23276 2596 23304
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 4430 23304 4436 23316
rect 4391 23276 4436 23304
rect 4430 23264 4436 23276
rect 4488 23264 4494 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 7101 23307 7159 23313
rect 7101 23304 7113 23307
rect 5960 23276 7113 23304
rect 5960 23264 5966 23276
rect 7101 23273 7113 23276
rect 7147 23304 7159 23307
rect 8110 23304 8116 23316
rect 7147 23276 8116 23304
rect 7147 23273 7159 23276
rect 7101 23267 7159 23273
rect 8110 23264 8116 23276
rect 8168 23264 8174 23316
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 11572 23276 11621 23304
rect 11572 23264 11578 23276
rect 11609 23273 11621 23276
rect 11655 23273 11667 23307
rect 12250 23304 12256 23316
rect 12211 23276 12256 23304
rect 11609 23267 11667 23273
rect 4982 23236 4988 23248
rect 4943 23208 4988 23236
rect 4982 23196 4988 23208
rect 5040 23196 5046 23248
rect 5718 23196 5724 23248
rect 5776 23196 5782 23248
rect 6362 23196 6368 23248
rect 6420 23236 6426 23248
rect 6733 23239 6791 23245
rect 6733 23236 6745 23239
rect 6420 23208 6745 23236
rect 6420 23196 6426 23208
rect 6733 23205 6745 23208
rect 6779 23205 6791 23239
rect 6733 23199 6791 23205
rect 1578 23168 1584 23180
rect 1539 23140 1584 23168
rect 1578 23128 1584 23140
rect 1636 23168 1642 23180
rect 1854 23168 1860 23180
rect 1636 23140 1860 23168
rect 1636 23128 1642 23140
rect 1854 23128 1860 23140
rect 1912 23128 1918 23180
rect 7190 23128 7196 23180
rect 7248 23168 7254 23180
rect 7561 23171 7619 23177
rect 7561 23168 7573 23171
rect 7248 23140 7573 23168
rect 7248 23128 7254 23140
rect 7561 23137 7573 23140
rect 7607 23168 7619 23171
rect 8294 23168 8300 23180
rect 7607 23140 8300 23168
rect 7607 23137 7619 23140
rect 7561 23131 7619 23137
rect 8294 23128 8300 23140
rect 8352 23128 8358 23180
rect 8570 23168 8576 23180
rect 8531 23140 8576 23168
rect 8570 23128 8576 23140
rect 8628 23128 8634 23180
rect 9309 23171 9367 23177
rect 9309 23137 9321 23171
rect 9355 23168 9367 23171
rect 9858 23168 9864 23180
rect 9355 23140 9864 23168
rect 9355 23137 9367 23140
rect 9309 23131 9367 23137
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 11624 23168 11652 23267
rect 12250 23264 12256 23276
rect 12308 23264 12314 23316
rect 12802 23264 12808 23316
rect 12860 23304 12866 23316
rect 13817 23307 13875 23313
rect 13817 23304 13829 23307
rect 12860 23276 13829 23304
rect 12860 23264 12866 23276
rect 13817 23273 13829 23276
rect 13863 23273 13875 23307
rect 13817 23267 13875 23273
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 16390 23304 16396 23316
rect 15611 23276 16396 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 18506 23304 18512 23316
rect 18467 23276 18512 23304
rect 18506 23264 18512 23276
rect 18564 23264 18570 23316
rect 19150 23304 19156 23316
rect 19111 23276 19156 23304
rect 19150 23264 19156 23276
rect 19208 23264 19214 23316
rect 19978 23304 19984 23316
rect 19939 23276 19984 23304
rect 19978 23264 19984 23276
rect 20036 23264 20042 23316
rect 16758 23196 16764 23248
rect 16816 23196 16822 23248
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19334 23236 19340 23248
rect 18923 23208 19340 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19334 23196 19340 23208
rect 19392 23236 19398 23248
rect 19613 23239 19671 23245
rect 19613 23236 19625 23239
rect 19392 23208 19625 23236
rect 19392 23196 19398 23208
rect 19613 23205 19625 23208
rect 19659 23236 19671 23239
rect 20162 23236 20168 23248
rect 19659 23208 20168 23236
rect 19659 23205 19671 23208
rect 19613 23199 19671 23205
rect 20162 23196 20168 23208
rect 20220 23236 20226 23248
rect 21174 23236 21180 23248
rect 20220 23208 21180 23236
rect 20220 23196 20226 23208
rect 21174 23196 21180 23208
rect 21232 23196 21238 23248
rect 11624 23140 12572 23168
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2866 23100 2872 23112
rect 2271 23072 2872 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 4709 23103 4767 23109
rect 4709 23100 4721 23103
rect 4126 23072 4721 23100
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 1765 22967 1823 22973
rect 1765 22964 1777 22967
rect 1728 22936 1777 22964
rect 1728 22924 1734 22936
rect 1765 22933 1777 22936
rect 1811 22933 1823 22967
rect 1765 22927 1823 22933
rect 2130 22924 2136 22976
rect 2188 22964 2194 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2188 22936 2973 22964
rect 2188 22924 2194 22936
rect 2961 22933 2973 22936
rect 3007 22964 3019 22967
rect 3602 22964 3608 22976
rect 3007 22936 3608 22964
rect 3007 22933 3019 22936
rect 2961 22927 3019 22933
rect 3602 22924 3608 22936
rect 3660 22964 3666 22976
rect 4126 22964 4154 23072
rect 4709 23069 4721 23072
rect 4755 23069 4767 23103
rect 12434 23100 12440 23112
rect 12395 23072 12440 23100
rect 4709 23063 4767 23069
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 12544 23100 12572 23140
rect 12618 23128 12624 23180
rect 12676 23168 12682 23180
rect 12989 23171 13047 23177
rect 12676 23140 12721 23168
rect 12676 23128 12682 23140
rect 12989 23137 13001 23171
rect 13035 23168 13047 23171
rect 13538 23168 13544 23180
rect 13035 23140 13544 23168
rect 13035 23137 13047 23140
rect 12989 23131 13047 23137
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 23014 23168 23020 23180
rect 22975 23140 23020 23168
rect 23014 23128 23020 23140
rect 23072 23128 23078 23180
rect 12897 23103 12955 23109
rect 12897 23100 12909 23103
rect 12544 23072 12909 23100
rect 12897 23069 12909 23072
rect 12943 23100 12955 23103
rect 13446 23100 13452 23112
rect 12943 23072 13452 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 15930 23100 15936 23112
rect 14323 23072 15936 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 16206 23100 16212 23112
rect 16167 23072 16212 23100
rect 16206 23060 16212 23072
rect 16264 23060 16270 23112
rect 16574 23060 16580 23112
rect 16632 23100 16638 23112
rect 17957 23103 18015 23109
rect 17957 23100 17969 23103
rect 16632 23072 17969 23100
rect 16632 23060 16638 23072
rect 17957 23069 17969 23072
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23100 21511 23103
rect 22002 23100 22008 23112
rect 21499 23072 22008 23100
rect 21499 23069 21511 23072
rect 21453 23063 21511 23069
rect 22002 23060 22008 23072
rect 22060 23060 22066 23112
rect 22830 23100 22836 23112
rect 22791 23072 22836 23100
rect 22830 23060 22836 23072
rect 22888 23060 22894 23112
rect 10781 23035 10839 23041
rect 10781 23001 10793 23035
rect 10827 23032 10839 23035
rect 11238 23032 11244 23044
rect 10827 23004 11244 23032
rect 10827 23001 10839 23004
rect 10781 22995 10839 23001
rect 11238 22992 11244 23004
rect 11296 22992 11302 23044
rect 12452 23032 12480 23060
rect 14642 23032 14648 23044
rect 12452 23004 14648 23032
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 21542 22992 21548 23044
rect 21600 23032 21606 23044
rect 22097 23035 22155 23041
rect 22097 23032 22109 23035
rect 21600 23004 22109 23032
rect 21600 22992 21606 23004
rect 22097 23001 22109 23004
rect 22143 23001 22155 23035
rect 22097 22995 22155 23001
rect 3660 22936 4154 22964
rect 3660 22924 3666 22936
rect 6086 22924 6092 22976
rect 6144 22964 6150 22976
rect 7745 22967 7803 22973
rect 7745 22964 7757 22967
rect 6144 22936 7757 22964
rect 6144 22924 6150 22936
rect 7745 22933 7757 22936
rect 7791 22933 7803 22967
rect 7745 22927 7803 22933
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 8757 22967 8815 22973
rect 8757 22964 8769 22967
rect 8260 22936 8769 22964
rect 8260 22924 8266 22936
rect 8757 22933 8769 22936
rect 8803 22933 8815 22967
rect 8757 22927 8815 22933
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10045 22967 10103 22973
rect 10045 22964 10057 22967
rect 10008 22936 10057 22964
rect 10008 22924 10014 22936
rect 10045 22933 10057 22936
rect 10091 22933 10103 22967
rect 10045 22927 10103 22933
rect 10413 22967 10471 22973
rect 10413 22933 10425 22967
rect 10459 22964 10471 22967
rect 10502 22964 10508 22976
rect 10459 22936 10508 22964
rect 10459 22933 10471 22936
rect 10413 22927 10471 22933
rect 10502 22924 10508 22936
rect 10560 22924 10566 22976
rect 10962 22924 10968 22976
rect 11020 22964 11026 22976
rect 11057 22967 11115 22973
rect 11057 22964 11069 22967
rect 11020 22936 11069 22964
rect 11020 22924 11026 22936
rect 11057 22933 11069 22936
rect 11103 22933 11115 22967
rect 11057 22927 11115 22933
rect 14921 22967 14979 22973
rect 14921 22933 14933 22967
rect 14967 22964 14979 22967
rect 15010 22964 15016 22976
rect 14967 22936 15016 22964
rect 14967 22933 14979 22936
rect 14921 22927 14979 22933
rect 15010 22924 15016 22936
rect 15068 22924 15074 22976
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21729 22967 21787 22973
rect 21729 22964 21741 22967
rect 21232 22936 21741 22964
rect 21232 22924 21238 22936
rect 21729 22933 21741 22936
rect 21775 22964 21787 22967
rect 22554 22964 22560 22976
rect 21775 22936 22560 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 1104 22874 24656 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 24656 22874
rect 1104 22800 24656 22822
rect 4801 22763 4859 22769
rect 4801 22729 4813 22763
rect 4847 22760 4859 22763
rect 4982 22760 4988 22772
rect 4847 22732 4988 22760
rect 4847 22729 4859 22732
rect 4801 22723 4859 22729
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 5169 22763 5227 22769
rect 5169 22729 5181 22763
rect 5215 22760 5227 22763
rect 5718 22760 5724 22772
rect 5215 22732 5724 22760
rect 5215 22729 5227 22732
rect 5169 22723 5227 22729
rect 5718 22720 5724 22732
rect 5776 22720 5782 22772
rect 7190 22760 7196 22772
rect 7151 22732 7196 22760
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 10870 22720 10876 22772
rect 10928 22760 10934 22772
rect 11977 22763 12035 22769
rect 11977 22760 11989 22763
rect 10928 22732 11989 22760
rect 10928 22720 10934 22732
rect 11977 22729 11989 22732
rect 12023 22760 12035 22763
rect 12434 22760 12440 22772
rect 12023 22732 12440 22760
rect 12023 22729 12035 22732
rect 11977 22723 12035 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 15841 22763 15899 22769
rect 15841 22729 15853 22763
rect 15887 22760 15899 22763
rect 16206 22760 16212 22772
rect 15887 22732 16212 22760
rect 15887 22729 15899 22732
rect 15841 22723 15899 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 18506 22720 18512 22772
rect 18564 22720 18570 22772
rect 23014 22760 23020 22772
rect 22975 22732 23020 22760
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 10502 22652 10508 22704
rect 10560 22692 10566 22704
rect 13170 22692 13176 22704
rect 10560 22664 11192 22692
rect 13131 22664 13176 22692
rect 10560 22652 10566 22664
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22624 1915 22627
rect 2406 22624 2412 22636
rect 1903 22596 2412 22624
rect 1903 22593 1915 22596
rect 1857 22587 1915 22593
rect 2406 22584 2412 22596
rect 2464 22584 2470 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10410 22624 10416 22636
rect 9999 22596 10416 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10410 22584 10416 22596
rect 10468 22624 10474 22636
rect 11164 22633 11192 22664
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 10468 22596 10701 22624
rect 10468 22584 10474 22596
rect 10689 22593 10701 22596
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22593 11207 22627
rect 14918 22624 14924 22636
rect 11149 22587 11207 22593
rect 13188 22596 14924 22624
rect 2130 22556 2136 22568
rect 2091 22528 2136 22556
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 5537 22559 5595 22565
rect 5537 22525 5549 22559
rect 5583 22525 5595 22559
rect 5537 22519 5595 22525
rect 7929 22559 7987 22565
rect 7929 22525 7941 22559
rect 7975 22525 7987 22559
rect 8386 22556 8392 22568
rect 8299 22528 8392 22556
rect 7929 22519 7987 22525
rect 2866 22448 2872 22500
rect 2924 22448 2930 22500
rect 4154 22448 4160 22500
rect 4212 22488 4218 22500
rect 4212 22460 4257 22488
rect 4212 22448 4218 22460
rect 4614 22380 4620 22432
rect 4672 22420 4678 22432
rect 5552 22420 5580 22519
rect 7944 22432 7972 22519
rect 8386 22516 8392 22528
rect 8444 22556 8450 22568
rect 10873 22559 10931 22565
rect 8444 22528 10272 22556
rect 8444 22516 8450 22528
rect 10244 22500 10272 22528
rect 10873 22525 10885 22559
rect 10919 22556 10931 22559
rect 10962 22556 10968 22568
rect 10919 22528 10968 22556
rect 10919 22525 10931 22528
rect 10873 22519 10931 22525
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 11238 22556 11244 22568
rect 11199 22528 11244 22556
rect 11238 22516 11244 22528
rect 11296 22516 11302 22568
rect 8478 22448 8484 22500
rect 8536 22448 8542 22500
rect 10226 22488 10232 22500
rect 10187 22460 10232 22488
rect 10226 22448 10232 22460
rect 10284 22448 10290 22500
rect 12989 22491 13047 22497
rect 12989 22457 13001 22491
rect 13035 22488 13047 22491
rect 13188 22488 13216 22596
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 15010 22584 15016 22636
rect 15068 22624 15074 22636
rect 16022 22624 16028 22636
rect 15068 22596 16028 22624
rect 15068 22584 15074 22596
rect 16022 22584 16028 22596
rect 16080 22624 16086 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16080 22596 16129 22624
rect 16080 22584 16086 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 18524 22624 18552 22720
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18524 22596 18705 22624
rect 16117 22587 16175 22593
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 20438 22624 20444 22636
rect 20399 22596 20444 22624
rect 18693 22587 18751 22593
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 16298 22556 16304 22568
rect 16259 22528 16304 22556
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 17313 22559 17371 22565
rect 17313 22525 17325 22559
rect 17359 22556 17371 22559
rect 17862 22556 17868 22568
rect 17359 22528 17868 22556
rect 17359 22525 17371 22528
rect 17313 22519 17371 22525
rect 17862 22516 17868 22528
rect 17920 22556 17926 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 17920 22528 18429 22556
rect 17920 22516 17926 22528
rect 18417 22525 18429 22528
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 21174 22516 21180 22568
rect 21232 22556 21238 22568
rect 21361 22559 21419 22565
rect 21361 22556 21373 22559
rect 21232 22528 21373 22556
rect 21232 22516 21238 22528
rect 21361 22525 21373 22528
rect 21407 22525 21419 22559
rect 21542 22556 21548 22568
rect 21503 22528 21548 22556
rect 21361 22519 21419 22525
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 22002 22516 22008 22568
rect 22060 22556 22066 22568
rect 22097 22559 22155 22565
rect 22097 22556 22109 22559
rect 22060 22528 22109 22556
rect 22060 22516 22066 22528
rect 22097 22525 22109 22528
rect 22143 22525 22155 22559
rect 22097 22519 22155 22525
rect 22281 22559 22339 22565
rect 22281 22525 22293 22559
rect 22327 22556 22339 22559
rect 22830 22556 22836 22568
rect 22327 22528 22836 22556
rect 22327 22525 22339 22528
rect 22281 22519 22339 22525
rect 13541 22491 13599 22497
rect 13541 22488 13553 22491
rect 13035 22460 13553 22488
rect 13035 22457 13047 22460
rect 12989 22451 13047 22457
rect 13541 22457 13553 22460
rect 13587 22457 13599 22491
rect 13541 22451 13599 22457
rect 13998 22448 14004 22500
rect 14056 22448 14062 22500
rect 15286 22488 15292 22500
rect 15247 22460 15292 22488
rect 15286 22448 15292 22460
rect 15344 22448 15350 22500
rect 18046 22488 18052 22500
rect 15580 22460 18052 22488
rect 5997 22423 6055 22429
rect 5997 22420 6009 22423
rect 4672 22392 6009 22420
rect 4672 22380 4678 22392
rect 5997 22389 6009 22392
rect 6043 22389 6055 22423
rect 5997 22383 6055 22389
rect 6178 22380 6184 22432
rect 6236 22420 6242 22432
rect 6365 22423 6423 22429
rect 6365 22420 6377 22423
rect 6236 22392 6377 22420
rect 6236 22380 6242 22392
rect 6365 22389 6377 22392
rect 6411 22389 6423 22423
rect 7926 22420 7932 22432
rect 7839 22392 7932 22420
rect 6365 22383 6423 22389
rect 7926 22380 7932 22392
rect 7984 22420 7990 22432
rect 8846 22420 8852 22432
rect 7984 22392 8852 22420
rect 7984 22380 7990 22392
rect 8846 22380 8852 22392
rect 8904 22420 8910 22432
rect 9950 22420 9956 22432
rect 8904 22392 9956 22420
rect 8904 22380 8910 22392
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 10870 22380 10876 22432
rect 10928 22420 10934 22432
rect 15580 22420 15608 22460
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 19150 22448 19156 22500
rect 19208 22448 19214 22500
rect 21085 22491 21143 22497
rect 21085 22457 21097 22491
rect 21131 22488 21143 22491
rect 22296 22488 22324 22519
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 21131 22460 22324 22488
rect 21131 22457 21143 22460
rect 21085 22451 21143 22457
rect 10928 22392 15608 22420
rect 17681 22423 17739 22429
rect 10928 22380 10934 22392
rect 17681 22389 17693 22423
rect 17727 22420 17739 22423
rect 19168 22420 19196 22448
rect 17727 22392 19196 22420
rect 17727 22389 17739 22392
rect 17681 22383 17739 22389
rect 21818 22380 21824 22432
rect 21876 22420 21882 22432
rect 22557 22423 22615 22429
rect 22557 22420 22569 22423
rect 21876 22392 22569 22420
rect 21876 22380 21882 22392
rect 22557 22389 22569 22392
rect 22603 22389 22615 22423
rect 22557 22383 22615 22389
rect 1104 22330 24656 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 24656 22330
rect 1104 22256 24656 22278
rect 1578 22216 1584 22228
rect 1539 22188 1584 22216
rect 1578 22176 1584 22188
rect 1636 22176 1642 22228
rect 3513 22219 3571 22225
rect 3513 22185 3525 22219
rect 3559 22216 3571 22219
rect 4154 22216 4160 22228
rect 3559 22188 4160 22216
rect 3559 22185 3571 22188
rect 3513 22179 3571 22185
rect 2590 22040 2596 22092
rect 2648 22080 2654 22092
rect 3053 22083 3111 22089
rect 3053 22080 3065 22083
rect 2648 22052 3065 22080
rect 2648 22040 2654 22052
rect 3053 22049 3065 22052
rect 3099 22080 3111 22083
rect 3528 22080 3556 22179
rect 4154 22176 4160 22188
rect 4212 22216 4218 22228
rect 4249 22219 4307 22225
rect 4249 22216 4261 22219
rect 4212 22188 4261 22216
rect 4212 22176 4218 22188
rect 4249 22185 4261 22188
rect 4295 22185 4307 22219
rect 4249 22179 4307 22185
rect 7561 22219 7619 22225
rect 7561 22185 7573 22219
rect 7607 22216 7619 22219
rect 7926 22216 7932 22228
rect 7607 22188 7932 22216
rect 7607 22185 7619 22188
rect 7561 22179 7619 22185
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 8570 22216 8576 22228
rect 8531 22188 8576 22216
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 11606 22216 11612 22228
rect 11567 22188 11612 22216
rect 11606 22176 11612 22188
rect 11664 22176 11670 22228
rect 13357 22219 13415 22225
rect 13357 22185 13369 22219
rect 13403 22216 13415 22219
rect 13998 22216 14004 22228
rect 13403 22188 14004 22216
rect 13403 22185 13415 22188
rect 13357 22179 13415 22185
rect 13998 22176 14004 22188
rect 14056 22216 14062 22228
rect 14369 22219 14427 22225
rect 14369 22216 14381 22219
rect 14056 22188 14381 22216
rect 14056 22176 14062 22188
rect 14369 22185 14381 22188
rect 14415 22185 14427 22219
rect 14369 22179 14427 22185
rect 14737 22219 14795 22225
rect 14737 22185 14749 22219
rect 14783 22216 14795 22219
rect 15286 22216 15292 22228
rect 14783 22188 15292 22216
rect 14783 22185 14795 22188
rect 14737 22179 14795 22185
rect 5718 22108 5724 22160
rect 5776 22108 5782 22160
rect 9309 22151 9367 22157
rect 9309 22117 9321 22151
rect 9355 22148 9367 22151
rect 11238 22148 11244 22160
rect 9355 22120 11244 22148
rect 9355 22117 9367 22120
rect 9309 22111 9367 22117
rect 5350 22080 5356 22092
rect 3099 22052 3556 22080
rect 5311 22052 5356 22080
rect 3099 22049 3111 22052
rect 3053 22043 3111 22049
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 6086 22080 6092 22092
rect 6047 22052 6092 22080
rect 6086 22040 6092 22052
rect 6144 22040 6150 22092
rect 7929 22083 7987 22089
rect 7929 22049 7941 22083
rect 7975 22080 7987 22083
rect 8386 22080 8392 22092
rect 7975 22052 8392 22080
rect 7975 22049 7987 22052
rect 7929 22043 7987 22049
rect 8386 22040 8392 22052
rect 8444 22040 8450 22092
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22080 10103 22083
rect 10226 22080 10232 22092
rect 10091 22052 10232 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 10502 22080 10508 22092
rect 10463 22052 10508 22080
rect 10502 22040 10508 22052
rect 10560 22040 10566 22092
rect 10612 22089 10640 22120
rect 11238 22108 11244 22120
rect 11296 22148 11302 22160
rect 11885 22151 11943 22157
rect 11885 22148 11897 22151
rect 11296 22120 11897 22148
rect 11296 22108 11302 22120
rect 11885 22117 11897 22120
rect 11931 22117 11943 22151
rect 11885 22111 11943 22117
rect 12618 22108 12624 22160
rect 12676 22148 12682 22160
rect 14752 22148 14780 22179
rect 15286 22176 15292 22188
rect 15344 22176 15350 22228
rect 16025 22219 16083 22225
rect 16025 22185 16037 22219
rect 16071 22216 16083 22219
rect 16758 22216 16764 22228
rect 16071 22188 16764 22216
rect 16071 22185 16083 22188
rect 16025 22179 16083 22185
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 12676 22120 14780 22148
rect 12676 22108 12682 22120
rect 18598 22108 18604 22160
rect 18656 22108 18662 22160
rect 19889 22151 19947 22157
rect 19889 22117 19901 22151
rect 19935 22148 19947 22151
rect 19978 22148 19984 22160
rect 19935 22120 19984 22148
rect 19935 22117 19947 22120
rect 19889 22111 19947 22117
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 20533 22151 20591 22157
rect 20533 22117 20545 22151
rect 20579 22148 20591 22151
rect 20579 22120 21588 22148
rect 20579 22117 20591 22120
rect 20533 22111 20591 22117
rect 21560 22092 21588 22120
rect 22094 22108 22100 22160
rect 22152 22108 22158 22160
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 10962 22040 10968 22092
rect 11020 22080 11026 22092
rect 12529 22083 12587 22089
rect 12529 22080 12541 22083
rect 11020 22052 12541 22080
rect 11020 22040 11026 22052
rect 12529 22049 12541 22052
rect 12575 22080 12587 22083
rect 12986 22080 12992 22092
rect 12575 22052 12992 22080
rect 12575 22049 12587 22052
rect 12529 22043 12587 22049
rect 12986 22040 12992 22052
rect 13044 22040 13050 22092
rect 14182 22080 14188 22092
rect 14143 22052 14188 22080
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 16574 22080 16580 22092
rect 16535 22052 16580 22080
rect 16574 22040 16580 22052
rect 16632 22040 16638 22092
rect 17589 22083 17647 22089
rect 17589 22049 17601 22083
rect 17635 22080 17647 22083
rect 17862 22080 17868 22092
rect 17635 22052 17868 22080
rect 17635 22049 17647 22052
rect 17589 22043 17647 22049
rect 2314 21972 2320 22024
rect 2372 22012 2378 22024
rect 2409 22015 2467 22021
rect 2409 22012 2421 22015
rect 2372 21984 2421 22012
rect 2372 21972 2378 21984
rect 2409 21981 2421 21984
rect 2455 21981 2467 22015
rect 9950 22012 9956 22024
rect 9911 21984 9956 22012
rect 2409 21975 2467 21981
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 12897 22015 12955 22021
rect 12897 22012 12909 22015
rect 12676 21984 12909 22012
rect 12676 21972 12682 21984
rect 12897 21981 12909 21984
rect 12943 22012 12955 22015
rect 13170 22012 13176 22024
rect 12943 21984 13176 22012
rect 12943 21981 12955 21984
rect 12897 21975 12955 21981
rect 13170 21972 13176 21984
rect 13228 22012 13234 22024
rect 13725 22015 13783 22021
rect 13725 22012 13737 22015
rect 13228 21984 13737 22012
rect 13228 21972 13234 21984
rect 13725 21981 13737 21984
rect 13771 22012 13783 22015
rect 14734 22012 14740 22024
rect 13771 21984 14740 22012
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 14734 21972 14740 21984
rect 14792 22012 14798 22024
rect 15657 22015 15715 22021
rect 15657 22012 15669 22015
rect 14792 21984 15669 22012
rect 14792 21972 14798 21984
rect 15657 21981 15669 21984
rect 15703 22012 15715 22015
rect 15930 22012 15936 22024
rect 15703 21984 15936 22012
rect 15703 21981 15715 21984
rect 15657 21975 15715 21981
rect 15930 21972 15936 21984
rect 15988 22012 15994 22024
rect 17604 22012 17632 22043
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 21174 22080 21180 22092
rect 21135 22052 21180 22080
rect 21174 22040 21180 22052
rect 21232 22040 21238 22092
rect 21542 22040 21548 22092
rect 21600 22080 21606 22092
rect 21729 22083 21787 22089
rect 21729 22080 21741 22083
rect 21600 22052 21741 22080
rect 21600 22040 21606 22052
rect 21729 22049 21741 22052
rect 21775 22049 21787 22083
rect 21729 22043 21787 22049
rect 18138 22012 18144 22024
rect 15988 21984 17632 22012
rect 18099 21984 18144 22012
rect 15988 21972 15994 21984
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 10965 21947 11023 21953
rect 10965 21944 10977 21947
rect 9732 21916 10977 21944
rect 9732 21904 9738 21916
rect 10965 21913 10977 21916
rect 11011 21913 11023 21947
rect 10965 21907 11023 21913
rect 2041 21879 2099 21885
rect 2041 21845 2053 21879
rect 2087 21876 2099 21879
rect 2498 21876 2504 21888
rect 2087 21848 2504 21876
rect 2087 21845 2099 21848
rect 2041 21839 2099 21845
rect 2498 21836 2504 21848
rect 2556 21836 2562 21888
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 23293 21879 23351 21885
rect 23293 21876 23305 21879
rect 22244 21848 23305 21876
rect 22244 21836 22250 21848
rect 23293 21845 23305 21848
rect 23339 21845 23351 21879
rect 23293 21839 23351 21845
rect 1104 21786 24656 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 24656 21786
rect 1104 21712 24656 21734
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 4157 21675 4215 21681
rect 4157 21672 4169 21675
rect 2924 21644 4169 21672
rect 2924 21632 2930 21644
rect 4157 21641 4169 21644
rect 4203 21641 4215 21675
rect 4157 21635 4215 21641
rect 5261 21675 5319 21681
rect 5261 21641 5273 21675
rect 5307 21672 5319 21675
rect 5350 21672 5356 21684
rect 5307 21644 5356 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 8386 21672 8392 21684
rect 8347 21644 8392 21672
rect 8386 21632 8392 21644
rect 8444 21632 8450 21684
rect 11974 21672 11980 21684
rect 11935 21644 11980 21672
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 16209 21675 16267 21681
rect 16209 21641 16221 21675
rect 16255 21672 16267 21675
rect 16298 21672 16304 21684
rect 16255 21644 16304 21672
rect 16255 21641 16267 21644
rect 16209 21635 16267 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 17681 21675 17739 21681
rect 17681 21641 17693 21675
rect 17727 21672 17739 21675
rect 18138 21672 18144 21684
rect 17727 21644 18144 21672
rect 17727 21641 17739 21644
rect 17681 21635 17739 21641
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22888 21644 23029 21672
rect 22888 21632 22894 21644
rect 23017 21641 23029 21644
rect 23063 21641 23075 21675
rect 23017 21635 23075 21641
rect 4893 21607 4951 21613
rect 4893 21573 4905 21607
rect 4939 21604 4951 21607
rect 5626 21604 5632 21616
rect 4939 21576 5632 21604
rect 4939 21573 4951 21576
rect 4893 21567 4951 21573
rect 5626 21564 5632 21576
rect 5684 21604 5690 21616
rect 6086 21604 6092 21616
rect 5684 21576 6092 21604
rect 5684 21564 5690 21576
rect 6086 21564 6092 21576
rect 6144 21564 6150 21616
rect 2498 21496 2504 21548
rect 2556 21536 2562 21548
rect 2869 21539 2927 21545
rect 2869 21536 2881 21539
rect 2556 21508 2881 21536
rect 2556 21496 2562 21508
rect 2869 21505 2881 21508
rect 2915 21505 2927 21539
rect 2869 21499 2927 21505
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21536 9183 21539
rect 9674 21536 9680 21548
rect 9171 21508 9680 21536
rect 9171 21505 9183 21508
rect 9125 21499 9183 21505
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 10410 21496 10416 21548
rect 10468 21536 10474 21548
rect 11425 21539 11483 21545
rect 11425 21536 11437 21539
rect 10468 21508 11437 21536
rect 10468 21496 10474 21508
rect 11425 21505 11437 21508
rect 11471 21505 11483 21539
rect 11992 21536 12020 21632
rect 17313 21607 17371 21613
rect 17313 21573 17325 21607
rect 17359 21604 17371 21607
rect 18598 21604 18604 21616
rect 17359 21576 18604 21604
rect 17359 21573 17371 21576
rect 17313 21567 17371 21573
rect 18598 21564 18604 21576
rect 18656 21604 18662 21616
rect 20257 21607 20315 21613
rect 20257 21604 20269 21607
rect 18656 21576 20269 21604
rect 18656 21564 18662 21576
rect 20257 21573 20269 21576
rect 20303 21573 20315 21607
rect 20257 21567 20315 21573
rect 21269 21607 21327 21613
rect 21269 21573 21281 21607
rect 21315 21604 21327 21607
rect 21315 21576 22324 21604
rect 21315 21573 21327 21576
rect 21269 21567 21327 21573
rect 12897 21539 12955 21545
rect 12897 21536 12909 21539
rect 11992 21508 12909 21536
rect 11425 21499 11483 21505
rect 12897 21505 12909 21508
rect 12943 21505 12955 21539
rect 12897 21499 12955 21505
rect 12986 21496 12992 21548
rect 13044 21536 13050 21548
rect 14645 21539 14703 21545
rect 14645 21536 14657 21539
rect 13044 21508 14657 21536
rect 13044 21496 13050 21508
rect 14645 21505 14657 21508
rect 14691 21505 14703 21539
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 14645 21499 14703 21505
rect 18984 21508 19165 21536
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 2130 21468 2136 21480
rect 1719 21440 2136 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 2130 21428 2136 21440
rect 2188 21468 2194 21480
rect 2409 21471 2467 21477
rect 2409 21468 2421 21471
rect 2188 21440 2421 21468
rect 2188 21428 2194 21440
rect 2409 21437 2421 21440
rect 2455 21437 2467 21471
rect 2590 21468 2596 21480
rect 2551 21440 2596 21468
rect 2409 21431 2467 21437
rect 2590 21428 2596 21440
rect 2648 21428 2654 21480
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 3973 21471 4031 21477
rect 3973 21437 3985 21471
rect 4019 21468 4031 21471
rect 4019 21440 4154 21468
rect 4019 21437 4031 21440
rect 3973 21431 4031 21437
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2976 21400 3004 21431
rect 3421 21403 3479 21409
rect 3421 21400 3433 21403
rect 2372 21372 3433 21400
rect 2372 21360 2378 21372
rect 3421 21369 3433 21372
rect 3467 21369 3479 21403
rect 3421 21363 3479 21369
rect 2222 21332 2228 21344
rect 2183 21304 2228 21332
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 4126 21332 4154 21440
rect 8570 21428 8576 21480
rect 8628 21468 8634 21480
rect 9401 21471 9459 21477
rect 9401 21468 9413 21471
rect 8628 21440 9413 21468
rect 8628 21428 8634 21440
rect 9401 21437 9413 21440
rect 9447 21437 9459 21471
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 9401 21431 9459 21437
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 18380 21440 18705 21468
rect 18380 21428 18386 21440
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18874 21468 18880 21480
rect 18835 21440 18880 21468
rect 18693 21431 18751 21437
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 8757 21403 8815 21409
rect 8757 21369 8769 21403
rect 8803 21400 8815 21403
rect 10134 21400 10140 21412
rect 8803 21372 10140 21400
rect 8803 21369 8815 21372
rect 8757 21363 8815 21369
rect 10134 21360 10140 21372
rect 10192 21360 10198 21412
rect 13354 21360 13360 21412
rect 13412 21360 13418 21412
rect 16942 21360 16948 21412
rect 17000 21400 17006 21412
rect 18233 21403 18291 21409
rect 18233 21400 18245 21403
rect 17000 21372 18245 21400
rect 17000 21360 17006 21372
rect 18233 21369 18245 21372
rect 18279 21369 18291 21403
rect 18233 21363 18291 21369
rect 18598 21360 18604 21412
rect 18656 21400 18662 21412
rect 18984 21400 19012 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 21542 21536 21548 21548
rect 21503 21508 21548 21536
rect 19153 21499 19211 21505
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 22296 21545 22324 21576
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21536 22339 21539
rect 23014 21536 23020 21548
rect 22327 21508 23020 21536
rect 22327 21505 22339 21508
rect 22281 21499 22339 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 19242 21468 19248 21480
rect 19203 21440 19248 21468
rect 19242 21428 19248 21440
rect 19300 21428 19306 21480
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21468 20131 21471
rect 22186 21468 22192 21480
rect 20119 21440 20668 21468
rect 22147 21440 22192 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 18656 21372 19012 21400
rect 19260 21400 19288 21428
rect 19705 21403 19763 21409
rect 19705 21400 19717 21403
rect 19260 21372 19717 21400
rect 18656 21360 18662 21372
rect 19705 21369 19717 21372
rect 19751 21369 19763 21403
rect 19705 21363 19763 21369
rect 4525 21335 4583 21341
rect 4525 21332 4537 21335
rect 4126 21304 4537 21332
rect 4525 21301 4537 21304
rect 4571 21332 4583 21335
rect 4614 21332 4620 21344
rect 4571 21304 4620 21332
rect 4571 21301 4583 21304
rect 4525 21295 4583 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 14918 21332 14924 21344
rect 14879 21304 14924 21332
rect 14918 21292 14924 21304
rect 14976 21332 14982 21344
rect 16574 21332 16580 21344
rect 14976 21304 16580 21332
rect 14976 21292 14982 21304
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 20640 21341 20668 21440
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 22554 21468 22560 21480
rect 22515 21440 22560 21468
rect 22554 21428 22560 21440
rect 22612 21428 22618 21480
rect 22741 21471 22799 21477
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 22830 21468 22836 21480
rect 22787 21440 22836 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 20625 21335 20683 21341
rect 20625 21301 20637 21335
rect 20671 21332 20683 21335
rect 21082 21332 21088 21344
rect 20671 21304 21088 21332
rect 20671 21301 20683 21304
rect 20625 21295 20683 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 1104 21242 24656 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 24656 21242
rect 1104 21168 24656 21190
rect 3602 21128 3608 21140
rect 3563 21100 3608 21128
rect 3602 21088 3608 21100
rect 3660 21088 3666 21140
rect 7834 21088 7840 21140
rect 7892 21128 7898 21140
rect 8570 21128 8576 21140
rect 7892 21100 8576 21128
rect 7892 21088 7898 21100
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 8846 21128 8852 21140
rect 8807 21100 8852 21128
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 12342 21128 12348 21140
rect 12303 21100 12348 21128
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 12713 21131 12771 21137
rect 12713 21097 12725 21131
rect 12759 21128 12771 21131
rect 13354 21128 13360 21140
rect 12759 21100 13360 21128
rect 12759 21097 12771 21100
rect 12713 21091 12771 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 14734 21128 14740 21140
rect 14695 21100 14740 21128
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 18322 21128 18328 21140
rect 18283 21100 18328 21128
rect 18322 21088 18328 21100
rect 18380 21088 18386 21140
rect 20533 21131 20591 21137
rect 20533 21097 20545 21131
rect 20579 21128 20591 21131
rect 21174 21128 21180 21140
rect 20579 21100 21180 21128
rect 20579 21097 20591 21100
rect 20533 21091 20591 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 21269 21131 21327 21137
rect 21269 21097 21281 21131
rect 21315 21128 21327 21131
rect 22002 21128 22008 21140
rect 21315 21100 22008 21128
rect 21315 21097 21327 21100
rect 21269 21091 21327 21097
rect 22002 21088 22008 21100
rect 22060 21128 22066 21140
rect 22554 21128 22560 21140
rect 22060 21100 22560 21128
rect 22060 21088 22066 21100
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 1670 21020 1676 21072
rect 1728 21060 1734 21072
rect 3237 21063 3295 21069
rect 3237 21060 3249 21063
rect 1728 21032 3249 21060
rect 1728 21020 1734 21032
rect 3237 21029 3249 21032
rect 3283 21029 3295 21063
rect 3237 21023 3295 21029
rect 5629 21063 5687 21069
rect 5629 21029 5641 21063
rect 5675 21060 5687 21063
rect 5718 21060 5724 21072
rect 5675 21032 5724 21060
rect 5675 21029 5687 21032
rect 5629 21023 5687 21029
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 6086 21020 6092 21072
rect 6144 21020 6150 21072
rect 7377 21063 7435 21069
rect 7377 21029 7389 21063
rect 7423 21060 7435 21063
rect 7650 21060 7656 21072
rect 7423 21032 7656 21060
rect 7423 21029 7435 21032
rect 7377 21023 7435 21029
rect 7650 21020 7656 21032
rect 7708 21020 7714 21072
rect 9309 21063 9367 21069
rect 9309 21029 9321 21063
rect 9355 21060 9367 21063
rect 9953 21063 10011 21069
rect 9953 21060 9965 21063
rect 9355 21032 9965 21060
rect 9355 21029 9367 21032
rect 9309 21023 9367 21029
rect 9953 21029 9965 21032
rect 9999 21060 10011 21063
rect 10502 21060 10508 21072
rect 9999 21032 10508 21060
rect 9999 21029 10011 21032
rect 9953 21023 10011 21029
rect 10502 21020 10508 21032
rect 10560 21020 10566 21072
rect 11885 21063 11943 21069
rect 11885 21029 11897 21063
rect 11931 21060 11943 21063
rect 12986 21060 12992 21072
rect 11931 21032 12992 21060
rect 11931 21029 11943 21032
rect 11885 21023 11943 21029
rect 12986 21020 12992 21032
rect 13044 21020 13050 21072
rect 17957 21063 18015 21069
rect 17957 21029 17969 21063
rect 18003 21060 18015 21063
rect 18138 21060 18144 21072
rect 18003 21032 18144 21060
rect 18003 21029 18015 21032
rect 17957 21023 18015 21029
rect 18138 21020 18144 21032
rect 18196 21020 18202 21072
rect 21818 21060 21824 21072
rect 21779 21032 21824 21060
rect 21818 21020 21824 21032
rect 21876 21020 21882 21072
rect 22370 21020 22376 21072
rect 22428 21020 22434 21072
rect 1765 20995 1823 21001
rect 1765 20961 1777 20995
rect 1811 20992 1823 20995
rect 2222 20992 2228 21004
rect 1811 20964 2228 20992
rect 1811 20961 1823 20964
rect 1765 20955 1823 20961
rect 2222 20952 2228 20964
rect 2280 20952 2286 21004
rect 2314 20952 2320 21004
rect 2372 20992 2378 21004
rect 2498 20992 2504 21004
rect 2372 20964 2417 20992
rect 2459 20964 2504 20992
rect 2372 20952 2378 20964
rect 2498 20952 2504 20964
rect 2556 20952 2562 21004
rect 4249 20995 4307 21001
rect 4249 20961 4261 20995
rect 4295 20992 4307 20995
rect 4614 20992 4620 21004
rect 4295 20964 4620 20992
rect 4295 20961 4307 20964
rect 4249 20955 4307 20961
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 10410 20992 10416 21004
rect 10371 20964 10416 20992
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 12161 20995 12219 21001
rect 12161 20992 12173 20995
rect 11480 20964 12173 20992
rect 11480 20952 11486 20964
rect 12161 20961 12173 20964
rect 12207 20961 12219 20995
rect 12161 20955 12219 20961
rect 13173 20995 13231 21001
rect 13173 20961 13185 20995
rect 13219 20992 13231 20995
rect 13814 20992 13820 21004
rect 13219 20964 13820 20992
rect 13219 20961 13231 20964
rect 13173 20955 13231 20961
rect 13814 20952 13820 20964
rect 13872 20992 13878 21004
rect 14182 20992 14188 21004
rect 13872 20964 14188 20992
rect 13872 20952 13878 20964
rect 14182 20952 14188 20964
rect 14240 20992 14246 21004
rect 14918 20992 14924 21004
rect 14240 20964 14924 20992
rect 14240 20952 14246 20964
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 16482 20992 16488 21004
rect 16443 20964 16488 20992
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 16942 20992 16948 21004
rect 16903 20964 16948 20992
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 18932 20964 19625 20992
rect 18932 20952 18938 20964
rect 19613 20961 19625 20964
rect 19659 20992 19671 20995
rect 20438 20992 20444 21004
rect 19659 20964 20444 20992
rect 19659 20961 19671 20964
rect 19613 20955 19671 20961
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 1670 20924 1676 20936
rect 1631 20896 1676 20924
rect 1670 20884 1676 20896
rect 1728 20884 1734 20936
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 6086 20924 6092 20936
rect 5399 20896 6092 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 2406 20816 2412 20868
rect 2464 20856 2470 20868
rect 2685 20859 2743 20865
rect 2685 20856 2697 20859
rect 2464 20828 2697 20856
rect 2464 20816 2470 20828
rect 2685 20825 2697 20828
rect 2731 20825 2743 20859
rect 2685 20819 2743 20825
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 4433 20859 4491 20865
rect 4433 20856 4445 20859
rect 3568 20828 4445 20856
rect 3568 20816 3574 20828
rect 4433 20825 4445 20828
rect 4479 20825 4491 20859
rect 4433 20819 4491 20825
rect 2038 20748 2044 20800
rect 2096 20788 2102 20800
rect 3602 20788 3608 20800
rect 2096 20760 3608 20788
rect 2096 20748 2102 20760
rect 3602 20748 3608 20760
rect 3660 20788 3666 20800
rect 5368 20788 5396 20887
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 18969 20927 19027 20933
rect 18969 20924 18981 20927
rect 17828 20896 18981 20924
rect 17828 20884 17834 20896
rect 18969 20893 18981 20896
rect 19015 20924 19027 20927
rect 19242 20924 19248 20936
rect 19015 20896 19248 20924
rect 19015 20893 19027 20896
rect 18969 20887 19027 20893
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20924 20131 20927
rect 21450 20924 21456 20936
rect 20119 20896 21456 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 7929 20859 7987 20865
rect 7929 20825 7941 20859
rect 7975 20856 7987 20859
rect 8570 20856 8576 20868
rect 7975 20828 8576 20856
rect 7975 20825 7987 20828
rect 7929 20819 7987 20825
rect 8570 20816 8576 20828
rect 8628 20816 8634 20868
rect 14369 20859 14427 20865
rect 14369 20825 14381 20859
rect 14415 20856 14427 20859
rect 14734 20856 14740 20868
rect 14415 20828 14740 20856
rect 14415 20825 14427 20828
rect 14369 20819 14427 20825
rect 14734 20816 14740 20828
rect 14792 20816 14798 20868
rect 19610 20816 19616 20868
rect 19668 20856 19674 20868
rect 20088 20856 20116 20887
rect 21450 20884 21456 20896
rect 21508 20924 21514 20936
rect 21545 20927 21603 20933
rect 21545 20924 21557 20927
rect 21508 20896 21557 20924
rect 21508 20884 21514 20896
rect 21545 20893 21557 20896
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 23014 20884 23020 20936
rect 23072 20924 23078 20936
rect 23569 20927 23627 20933
rect 23569 20924 23581 20927
rect 23072 20896 23581 20924
rect 23072 20884 23078 20896
rect 23569 20893 23581 20896
rect 23615 20893 23627 20927
rect 23569 20887 23627 20893
rect 19668 20828 20116 20856
rect 19668 20816 19674 20828
rect 18598 20788 18604 20800
rect 3660 20760 5396 20788
rect 18559 20760 18604 20788
rect 3660 20748 3666 20760
rect 18598 20748 18604 20760
rect 18656 20748 18662 20800
rect 1104 20698 24656 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 24656 20698
rect 1104 20624 24656 20646
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 5445 20587 5503 20593
rect 2188 20556 4200 20584
rect 2188 20544 2194 20556
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 2406 20448 2412 20460
rect 1903 20420 2412 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 4172 20457 4200 20556
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 5718 20584 5724 20596
rect 5491 20556 5724 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10192 20556 10885 20584
rect 10192 20544 10198 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 16393 20587 16451 20593
rect 16393 20553 16405 20587
rect 16439 20584 16451 20587
rect 16482 20584 16488 20596
rect 16439 20556 16488 20584
rect 16439 20553 16451 20556
rect 16393 20547 16451 20553
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 16761 20587 16819 20593
rect 16761 20553 16773 20587
rect 16807 20584 16819 20587
rect 16942 20584 16948 20596
rect 16807 20556 16948 20584
rect 16807 20553 16819 20556
rect 16761 20547 16819 20553
rect 16942 20544 16948 20556
rect 17000 20584 17006 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 17000 20556 17049 20584
rect 17000 20544 17006 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 17037 20547 17095 20553
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20584 18383 20587
rect 18874 20584 18880 20596
rect 18371 20556 18880 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 21913 20587 21971 20593
rect 21913 20584 21925 20587
rect 21876 20556 21925 20584
rect 21876 20544 21882 20556
rect 21913 20553 21925 20556
rect 21959 20553 21971 20587
rect 22370 20584 22376 20596
rect 22331 20556 22376 20584
rect 21913 20547 21971 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 10229 20519 10287 20525
rect 10229 20485 10241 20519
rect 10275 20516 10287 20519
rect 10410 20516 10416 20528
rect 10275 20488 10416 20516
rect 10275 20485 10287 20488
rect 10229 20479 10287 20485
rect 10410 20476 10416 20488
rect 10468 20476 10474 20528
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20417 4215 20451
rect 4157 20411 4215 20417
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 8113 20451 8171 20457
rect 8113 20448 8125 20451
rect 7607 20420 8125 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 8113 20417 8125 20420
rect 8159 20448 8171 20451
rect 8478 20448 8484 20460
rect 8159 20420 8484 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8478 20408 8484 20420
rect 8536 20408 8542 20460
rect 13998 20448 14004 20460
rect 13911 20420 14004 20448
rect 13998 20408 14004 20420
rect 14056 20448 14062 20460
rect 14642 20448 14648 20460
rect 14056 20420 14648 20448
rect 14056 20408 14062 20420
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20448 16083 20451
rect 16298 20448 16304 20460
rect 16071 20420 16304 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20448 19027 20451
rect 20346 20448 20352 20460
rect 19015 20420 20352 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 21637 20451 21695 20457
rect 21637 20448 21649 20451
rect 20496 20420 21649 20448
rect 20496 20408 20502 20420
rect 21637 20417 21649 20420
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2133 20383 2191 20389
rect 2133 20380 2145 20383
rect 2096 20352 2145 20380
rect 2096 20340 2102 20352
rect 2133 20349 2145 20352
rect 2179 20349 2191 20383
rect 2133 20343 2191 20349
rect 3510 20340 3516 20392
rect 3568 20340 3574 20392
rect 6086 20340 6092 20392
rect 6144 20380 6150 20392
rect 6181 20383 6239 20389
rect 6181 20380 6193 20383
rect 6144 20352 6193 20380
rect 6144 20340 6150 20352
rect 6181 20349 6193 20352
rect 6227 20380 6239 20383
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 6227 20352 7205 20380
rect 6227 20349 6239 20352
rect 6181 20343 6239 20349
rect 7193 20349 7205 20352
rect 7239 20380 7251 20383
rect 7834 20380 7840 20392
rect 7239 20352 7840 20380
rect 7239 20349 7251 20352
rect 7193 20343 7251 20349
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 10689 20383 10747 20389
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 13265 20383 13323 20389
rect 10735 20352 11284 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 8570 20272 8576 20324
rect 8628 20272 8634 20324
rect 9858 20312 9864 20324
rect 9819 20284 9864 20312
rect 9858 20272 9864 20284
rect 9916 20272 9922 20324
rect 4525 20247 4583 20253
rect 4525 20213 4537 20247
rect 4571 20244 4583 20247
rect 4614 20244 4620 20256
rect 4571 20216 4620 20244
rect 4571 20213 4583 20216
rect 4525 20207 4583 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5810 20244 5816 20256
rect 5771 20216 5816 20244
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 11256 20253 11284 20352
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 13722 20380 13728 20392
rect 13311 20352 13728 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 19610 20380 19616 20392
rect 19571 20352 19616 20380
rect 19610 20340 19616 20352
rect 19668 20340 19674 20392
rect 13633 20315 13691 20321
rect 13633 20281 13645 20315
rect 13679 20312 13691 20315
rect 14274 20312 14280 20324
rect 13679 20284 14280 20312
rect 13679 20281 13691 20284
rect 13633 20275 13691 20281
rect 14274 20272 14280 20284
rect 14332 20272 14338 20324
rect 14734 20272 14740 20324
rect 14792 20272 14798 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 19889 20315 19947 20321
rect 19889 20312 19901 20315
rect 19383 20284 19901 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 19889 20281 19901 20284
rect 19935 20281 19947 20315
rect 19889 20275 19947 20281
rect 11241 20247 11299 20253
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 11422 20244 11428 20256
rect 11287 20216 11428 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11422 20204 11428 20216
rect 11480 20204 11486 20256
rect 12713 20247 12771 20253
rect 12713 20213 12725 20247
rect 12759 20244 12771 20247
rect 12986 20244 12992 20256
rect 12759 20216 12992 20244
rect 12759 20213 12771 20216
rect 12713 20207 12771 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 13814 20244 13820 20256
rect 13780 20216 13820 20244
rect 13780 20204 13786 20216
rect 13814 20204 13820 20216
rect 13872 20244 13878 20256
rect 14458 20244 14464 20256
rect 13872 20216 14464 20244
rect 13872 20204 13878 20216
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 19904 20244 19932 20275
rect 20346 20272 20352 20324
rect 20404 20272 20410 20324
rect 22094 20244 22100 20256
rect 19904 20216 22100 20244
rect 22094 20204 22100 20216
rect 22152 20204 22158 20256
rect 1104 20154 24656 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 24656 20154
rect 1104 20080 24656 20102
rect 2133 20043 2191 20049
rect 2133 20009 2145 20043
rect 2179 20040 2191 20043
rect 3510 20040 3516 20052
rect 2179 20012 3516 20040
rect 2179 20009 2191 20012
rect 2133 20003 2191 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 14093 20043 14151 20049
rect 14093 20009 14105 20043
rect 14139 20040 14151 20043
rect 14734 20040 14740 20052
rect 14139 20012 14740 20040
rect 14139 20009 14151 20012
rect 14093 20003 14151 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 16669 20043 16727 20049
rect 16669 20040 16681 20043
rect 16540 20012 16681 20040
rect 16540 20000 16546 20012
rect 16669 20009 16681 20012
rect 16715 20009 16727 20043
rect 16669 20003 16727 20009
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19972 1731 19975
rect 2406 19972 2412 19984
rect 1719 19944 2412 19972
rect 1719 19941 1731 19944
rect 1673 19935 1731 19941
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 5813 19975 5871 19981
rect 5813 19941 5825 19975
rect 5859 19972 5871 19975
rect 6822 19972 6828 19984
rect 5859 19944 6828 19972
rect 5859 19941 5871 19944
rect 5813 19935 5871 19941
rect 6822 19932 6828 19944
rect 6880 19932 6886 19984
rect 2130 19864 2136 19916
rect 2188 19904 2194 19916
rect 2501 19907 2559 19913
rect 2501 19904 2513 19907
rect 2188 19876 2513 19904
rect 2188 19864 2194 19876
rect 2501 19873 2513 19876
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4798 19904 4804 19916
rect 4120 19876 4804 19904
rect 4120 19864 4126 19876
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 6086 19904 6092 19916
rect 6047 19876 6092 19904
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 9858 19904 9864 19916
rect 9364 19876 9864 19904
rect 9364 19864 9370 19876
rect 9858 19864 9864 19876
rect 9916 19904 9922 19916
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 9916 19876 9965 19904
rect 9916 19864 9922 19876
rect 9953 19873 9965 19876
rect 9999 19873 10011 19907
rect 11514 19904 11520 19916
rect 11475 19876 11520 19904
rect 9953 19867 10011 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19904 12955 19907
rect 12986 19904 12992 19916
rect 12943 19876 12992 19904
rect 12943 19873 12955 19876
rect 12897 19867 12955 19873
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 15930 19904 15936 19916
rect 15611 19876 15936 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 16684 19904 16712 20003
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 21269 20043 21327 20049
rect 21269 20040 21281 20043
rect 20404 20012 21281 20040
rect 20404 20000 20410 20012
rect 21269 20009 21281 20012
rect 21315 20009 21327 20043
rect 21269 20003 21327 20009
rect 16942 19932 16948 19984
rect 17000 19972 17006 19984
rect 18969 19975 19027 19981
rect 17000 19944 17264 19972
rect 17000 19932 17006 19944
rect 16758 19904 16764 19916
rect 16671 19876 16764 19904
rect 16758 19864 16764 19876
rect 16816 19904 16822 19916
rect 17236 19913 17264 19944
rect 18969 19941 18981 19975
rect 19015 19972 19027 19975
rect 20438 19972 20444 19984
rect 19015 19944 20444 19972
rect 19015 19941 19027 19944
rect 18969 19935 19027 19941
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 22554 19972 22560 19984
rect 22515 19944 22560 19972
rect 22554 19932 22560 19944
rect 22612 19932 22618 19984
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 16816 19876 17049 19904
rect 16816 19864 16822 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19873 17279 19907
rect 17770 19904 17776 19916
rect 17731 19876 17776 19904
rect 17221 19867 17279 19873
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 17954 19904 17960 19916
rect 17915 19876 17960 19904
rect 17954 19864 17960 19876
rect 18012 19904 18018 19916
rect 18012 19876 18276 19904
rect 18012 19864 18018 19876
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5718 19836 5724 19848
rect 5307 19808 5724 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 6362 19836 6368 19848
rect 6323 19808 6368 19836
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 8110 19836 8116 19848
rect 8071 19808 8116 19836
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 11146 19796 11152 19848
rect 11204 19836 11210 19848
rect 11333 19839 11391 19845
rect 11333 19836 11345 19839
rect 11204 19808 11345 19836
rect 11204 19796 11210 19808
rect 11333 19805 11345 19808
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 16022 19836 16028 19848
rect 15983 19808 16028 19836
rect 15473 19799 15531 19805
rect 15286 19728 15292 19780
rect 15344 19768 15350 19780
rect 15488 19768 15516 19799
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 18248 19836 18276 19876
rect 18322 19864 18328 19916
rect 18380 19904 18386 19916
rect 19337 19907 19395 19913
rect 19337 19904 19349 19907
rect 18380 19876 19349 19904
rect 18380 19864 18386 19876
rect 19337 19873 19349 19876
rect 19383 19904 19395 19907
rect 19426 19904 19432 19916
rect 19383 19876 19432 19904
rect 19383 19873 19395 19876
rect 19337 19867 19395 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 21082 19904 21088 19916
rect 21043 19876 21088 19904
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 22186 19864 22192 19916
rect 22244 19904 22250 19916
rect 22649 19907 22707 19913
rect 22649 19904 22661 19907
rect 22244 19876 22661 19904
rect 22244 19864 22250 19876
rect 22649 19873 22661 19876
rect 22695 19904 22707 19907
rect 22738 19904 22744 19916
rect 22695 19876 22744 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 18598 19836 18604 19848
rect 18248 19808 18604 19836
rect 18598 19796 18604 19808
rect 18656 19836 18662 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18656 19808 19257 19836
rect 18656 19796 18662 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 16114 19768 16120 19780
rect 15344 19740 16120 19768
rect 15344 19728 15350 19740
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 3510 19700 3516 19712
rect 3471 19672 3516 19700
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 9306 19700 9312 19712
rect 9267 19672 9312 19700
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 10318 19700 10324 19712
rect 10279 19672 10324 19700
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 13081 19703 13139 19709
rect 13081 19700 13093 19703
rect 12124 19672 13093 19700
rect 12124 19660 12130 19672
rect 13081 19669 13093 19672
rect 13127 19669 13139 19703
rect 14458 19700 14464 19712
rect 14419 19672 14464 19700
rect 13081 19663 13139 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 18233 19703 18291 19709
rect 18233 19669 18245 19703
rect 18279 19700 18291 19703
rect 18506 19700 18512 19712
rect 18279 19672 18512 19700
rect 18279 19669 18291 19672
rect 18233 19663 18291 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 21450 19660 21456 19712
rect 21508 19700 21514 19712
rect 21545 19703 21603 19709
rect 21545 19700 21557 19703
rect 21508 19672 21557 19700
rect 21508 19660 21514 19672
rect 21545 19669 21557 19672
rect 21591 19669 21603 19703
rect 21545 19663 21603 19669
rect 1104 19610 24656 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 24656 19610
rect 1104 19536 24656 19558
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 3789 19499 3847 19505
rect 3789 19496 3801 19499
rect 3568 19468 3801 19496
rect 3568 19456 3574 19468
rect 3789 19465 3801 19468
rect 3835 19465 3847 19499
rect 3789 19459 3847 19465
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 5350 19496 5356 19508
rect 5031 19468 5356 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5350 19456 5356 19468
rect 5408 19456 5414 19508
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 6362 19496 6368 19508
rect 6319 19468 6368 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8021 19499 8079 19505
rect 8021 19496 8033 19499
rect 7892 19468 8033 19496
rect 7892 19456 7898 19468
rect 8021 19465 8033 19468
rect 8067 19465 8079 19499
rect 8021 19459 8079 19465
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 9125 19499 9183 19505
rect 9125 19496 9137 19499
rect 8628 19468 9137 19496
rect 8628 19456 8634 19468
rect 9125 19465 9137 19468
rect 9171 19465 9183 19499
rect 16758 19496 16764 19508
rect 16719 19468 16764 19496
rect 9125 19459 9183 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 20901 19499 20959 19505
rect 20901 19496 20913 19499
rect 19116 19468 20913 19496
rect 19116 19456 19122 19468
rect 20901 19465 20913 19468
rect 20947 19496 20959 19499
rect 21082 19496 21088 19508
rect 20947 19468 21088 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22370 19496 22376 19508
rect 22143 19468 22376 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 22738 19496 22744 19508
rect 22699 19468 22744 19496
rect 22738 19456 22744 19468
rect 22796 19456 22802 19508
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19428 9735 19431
rect 9723 19400 10732 19428
rect 9723 19397 9735 19400
rect 9677 19391 9735 19397
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19360 4491 19363
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 4479 19332 5457 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 5445 19329 5457 19332
rect 5491 19360 5503 19363
rect 5491 19332 7144 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 7116 19304 7144 19332
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10704 19369 10732 19400
rect 10689 19363 10747 19369
rect 9916 19332 10640 19360
rect 9916 19320 9922 19332
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2222 19252 2228 19304
rect 2280 19292 2286 19304
rect 2501 19295 2559 19301
rect 2501 19292 2513 19295
rect 2280 19264 2513 19292
rect 2280 19252 2286 19264
rect 2501 19261 2513 19264
rect 2547 19292 2559 19295
rect 3510 19292 3516 19304
rect 2547 19264 3516 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19261 5411 19295
rect 5718 19292 5724 19304
rect 5679 19264 5724 19292
rect 5353 19255 5411 19261
rect 2406 19116 2412 19168
rect 2464 19156 2470 19168
rect 2608 19156 2636 19224
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 5368 19224 5396 19255
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19292 5963 19295
rect 6270 19292 6276 19304
rect 5951 19264 6276 19292
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 6270 19252 6276 19264
rect 6328 19292 6334 19304
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6328 19264 7021 19292
rect 6328 19252 6334 19264
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7156 19264 7665 19292
rect 7156 19252 7162 19264
rect 7653 19261 7665 19264
rect 7699 19292 7711 19295
rect 8110 19292 8116 19304
rect 7699 19264 8116 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 10612 19301 10640 19332
rect 10689 19329 10701 19363
rect 10735 19360 10747 19363
rect 11514 19360 11520 19372
rect 10735 19332 11520 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19360 17739 19363
rect 18506 19360 18512 19372
rect 17727 19332 18512 19360
rect 17727 19329 17739 19332
rect 17681 19323 17739 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 19576 19332 20269 19360
rect 19576 19320 19582 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 8665 19295 8723 19301
rect 8665 19261 8677 19295
rect 8711 19292 8723 19295
rect 8941 19295 8999 19301
rect 8941 19292 8953 19295
rect 8711 19264 8953 19292
rect 8711 19261 8723 19264
rect 8665 19255 8723 19261
rect 8941 19261 8953 19264
rect 8987 19292 8999 19295
rect 10597 19295 10655 19301
rect 8987 19264 10272 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 4120 19196 5396 19224
rect 4120 19184 4126 19196
rect 10042 19156 10048 19168
rect 2464 19128 2636 19156
rect 10003 19128 10048 19156
rect 2464 19116 2470 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10244 19156 10272 19264
rect 10597 19261 10609 19295
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19261 11023 19295
rect 11146 19292 11152 19304
rect 11107 19264 11152 19292
rect 10965 19255 11023 19261
rect 10318 19184 10324 19236
rect 10376 19224 10382 19236
rect 10980 19224 11008 19255
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 12069 19295 12127 19301
rect 12069 19261 12081 19295
rect 12115 19292 12127 19295
rect 12894 19292 12900 19304
rect 12115 19264 12900 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19292 13783 19295
rect 13998 19292 14004 19304
rect 13771 19264 14004 19292
rect 13771 19261 13783 19264
rect 13725 19255 13783 19261
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 14516 19264 15301 19292
rect 14516 19252 14522 19264
rect 15289 19261 15301 19264
rect 15335 19292 15347 19295
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 15335 19264 15577 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 11514 19224 11520 19236
rect 10376 19196 11008 19224
rect 11427 19196 11520 19224
rect 10376 19184 10382 19196
rect 11514 19184 11520 19196
rect 11572 19224 11578 19236
rect 12710 19224 12716 19236
rect 11572 19196 12716 19224
rect 11572 19184 11578 19196
rect 12710 19184 12716 19196
rect 12768 19184 12774 19236
rect 14274 19184 14280 19236
rect 14332 19184 14338 19236
rect 15580 19224 15608 19255
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 16574 19292 16580 19304
rect 16080 19264 16580 19292
rect 16080 19252 16086 19264
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 18230 19292 18236 19304
rect 18191 19264 18236 19292
rect 18230 19252 18236 19264
rect 18288 19252 18294 19304
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21913 19295 21971 19301
rect 21913 19292 21925 19295
rect 21140 19264 21925 19292
rect 21140 19252 21146 19264
rect 21913 19261 21925 19264
rect 21959 19292 21971 19295
rect 22278 19292 22284 19304
rect 21959 19264 22284 19292
rect 21959 19261 21971 19264
rect 21913 19255 21971 19261
rect 22278 19252 22284 19264
rect 22336 19292 22342 19304
rect 22373 19295 22431 19301
rect 22373 19292 22385 19295
rect 22336 19264 22385 19292
rect 22336 19252 22342 19264
rect 22373 19261 22385 19264
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 17310 19224 17316 19236
rect 15580 19196 17316 19224
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 19242 19184 19248 19236
rect 19300 19184 19306 19236
rect 11422 19156 11428 19168
rect 10244 19128 11428 19156
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 15746 19156 15752 19168
rect 15707 19128 15752 19156
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 16022 19156 16028 19168
rect 15983 19128 16028 19156
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 16172 19128 17141 19156
rect 16172 19116 16178 19128
rect 17129 19125 17141 19128
rect 17175 19156 17187 19159
rect 21726 19156 21732 19168
rect 17175 19128 21732 19156
rect 17175 19125 17187 19128
rect 17129 19119 17187 19125
rect 21726 19116 21732 19128
rect 21784 19116 21790 19168
rect 1104 19066 24656 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 24656 19066
rect 1104 18992 24656 19014
rect 1673 18955 1731 18961
rect 1673 18921 1685 18955
rect 1719 18952 1731 18955
rect 2314 18952 2320 18964
rect 1719 18924 2320 18952
rect 1719 18921 1731 18924
rect 1673 18915 1731 18921
rect 2314 18912 2320 18924
rect 2372 18912 2378 18964
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 5718 18952 5724 18964
rect 4479 18924 5724 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6362 18912 6368 18964
rect 6420 18952 6426 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 6420 18924 6561 18952
rect 6420 18912 6426 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 6549 18915 6607 18921
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 7745 18955 7803 18961
rect 7745 18952 7757 18955
rect 6880 18924 7757 18952
rect 6880 18912 6886 18924
rect 7745 18921 7757 18924
rect 7791 18921 7803 18955
rect 9306 18952 9312 18964
rect 9267 18924 9312 18952
rect 7745 18915 7803 18921
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10502 18952 10508 18964
rect 10091 18924 10508 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10502 18912 10508 18924
rect 10560 18952 10566 18964
rect 11146 18952 11152 18964
rect 10560 18924 11152 18952
rect 10560 18912 10566 18924
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14148 18924 14473 18952
rect 14148 18912 14154 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 16574 18952 16580 18964
rect 16535 18924 16580 18952
rect 14461 18915 14519 18921
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 17497 18955 17555 18961
rect 17497 18921 17509 18955
rect 17543 18952 17555 18955
rect 17770 18952 17776 18964
rect 17543 18924 17776 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 19242 18952 19248 18964
rect 18187 18924 19248 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19484 18924 19533 18952
rect 19484 18912 19490 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 2188 18856 2421 18884
rect 2188 18844 2194 18856
rect 2409 18853 2421 18856
rect 2455 18853 2467 18887
rect 2409 18847 2467 18853
rect 5350 18844 5356 18896
rect 5408 18844 5414 18896
rect 1670 18776 1676 18828
rect 1728 18816 1734 18828
rect 1949 18819 2007 18825
rect 1949 18816 1961 18819
rect 1728 18788 1961 18816
rect 1728 18776 1734 18788
rect 1949 18785 1961 18788
rect 1995 18785 2007 18819
rect 1949 18779 2007 18785
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 3050 18816 3056 18828
rect 3007 18788 3056 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 3050 18776 3056 18788
rect 3108 18816 3114 18828
rect 3108 18788 4154 18816
rect 3108 18776 3114 18788
rect 4126 18680 4154 18788
rect 5074 18776 5080 18828
rect 5132 18816 5138 18828
rect 5368 18816 5396 18844
rect 5491 18819 5549 18825
rect 5491 18816 5503 18819
rect 5132 18788 5503 18816
rect 5132 18776 5138 18788
rect 5491 18785 5503 18788
rect 5537 18785 5549 18819
rect 5736 18816 5764 18912
rect 7098 18884 7104 18896
rect 7059 18856 7104 18884
rect 7098 18844 7104 18856
rect 7156 18844 7162 18896
rect 12710 18884 12716 18896
rect 12671 18856 12716 18884
rect 12710 18844 12716 18856
rect 12768 18844 12774 18896
rect 17129 18887 17187 18893
rect 17129 18853 17141 18887
rect 17175 18884 17187 18887
rect 17954 18884 17960 18896
rect 17175 18856 17960 18884
rect 17175 18853 17187 18856
rect 17129 18847 17187 18853
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 21818 18844 21824 18896
rect 21876 18844 21882 18896
rect 22738 18844 22744 18896
rect 22796 18884 22802 18896
rect 23109 18887 23167 18893
rect 23109 18884 23121 18887
rect 22796 18856 23121 18884
rect 22796 18844 22802 18856
rect 23109 18853 23121 18856
rect 23155 18853 23167 18887
rect 23109 18847 23167 18853
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 5736 18788 6101 18816
rect 5491 18779 5549 18785
rect 6089 18785 6101 18788
rect 6135 18785 6147 18819
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6089 18779 6147 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 7834 18816 7840 18828
rect 7607 18788 7840 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 5350 18748 5356 18760
rect 5311 18720 5356 18748
rect 5350 18708 5356 18720
rect 5408 18748 5414 18760
rect 5626 18748 5632 18760
rect 5408 18720 5632 18748
rect 5408 18708 5414 18720
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 4614 18680 4620 18692
rect 4126 18652 4620 18680
rect 4614 18640 4620 18652
rect 4672 18680 4678 18692
rect 7576 18680 7604 18779
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 15930 18816 15936 18828
rect 15891 18788 15936 18816
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 19058 18816 19064 18828
rect 19019 18788 19064 18816
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10962 18748 10968 18760
rect 10923 18720 10968 18748
rect 10689 18711 10747 18717
rect 4672 18652 7604 18680
rect 4672 18640 4678 18652
rect 3142 18612 3148 18624
rect 3103 18584 3148 18612
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 4798 18612 4804 18624
rect 4759 18584 4804 18612
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 10318 18612 10324 18624
rect 10279 18584 10324 18612
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 10704 18612 10732 18711
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16390 18748 16396 18760
rect 16255 18720 16396 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20438 18748 20444 18760
rect 20027 18720 20444 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18717 21143 18751
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 21085 18711 21143 18717
rect 11054 18612 11060 18624
rect 10704 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 12986 18612 12992 18624
rect 11480 18584 12992 18612
rect 11480 18572 11486 18584
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13449 18615 13507 18621
rect 13449 18581 13461 18615
rect 13495 18612 13507 18615
rect 13998 18612 14004 18624
rect 13495 18584 14004 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18417 18615 18475 18621
rect 18417 18612 18429 18615
rect 18288 18584 18429 18612
rect 18288 18572 18294 18584
rect 18417 18581 18429 18584
rect 18463 18581 18475 18615
rect 18417 18575 18475 18581
rect 20533 18615 20591 18621
rect 20533 18581 20545 18615
rect 20579 18612 20591 18615
rect 21100 18612 21128 18711
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 21450 18612 21456 18624
rect 20579 18584 21456 18612
rect 20579 18581 20591 18584
rect 20533 18575 20591 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 24656 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 24656 18522
rect 1104 18448 24656 18470
rect 5074 18408 5080 18420
rect 5035 18380 5080 18408
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5718 18408 5724 18420
rect 5679 18380 5724 18408
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 7193 18411 7251 18417
rect 7193 18408 7205 18411
rect 5868 18380 7205 18408
rect 5868 18368 5874 18380
rect 7193 18377 7205 18380
rect 7239 18377 7251 18411
rect 7193 18371 7251 18377
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 10318 18408 10324 18420
rect 9263 18380 10324 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21453 18411 21511 18417
rect 21453 18408 21465 18411
rect 21416 18380 21465 18408
rect 21416 18368 21422 18380
rect 21453 18377 21465 18380
rect 21499 18408 21511 18411
rect 21729 18411 21787 18417
rect 21729 18408 21741 18411
rect 21499 18380 21741 18408
rect 21499 18377 21511 18380
rect 21453 18371 21511 18377
rect 21729 18377 21741 18380
rect 21775 18377 21787 18411
rect 21729 18371 21787 18377
rect 4798 18300 4804 18352
rect 4856 18340 4862 18352
rect 5445 18343 5503 18349
rect 5445 18340 5457 18343
rect 4856 18312 5457 18340
rect 4856 18300 4862 18312
rect 5445 18309 5457 18312
rect 5491 18340 5503 18343
rect 6270 18340 6276 18352
rect 5491 18312 6276 18340
rect 5491 18309 5503 18312
rect 5445 18303 5503 18309
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 10962 18340 10968 18352
rect 10923 18312 10968 18340
rect 10962 18300 10968 18312
rect 11020 18340 11026 18352
rect 11517 18343 11575 18349
rect 11517 18340 11529 18343
rect 11020 18312 11529 18340
rect 11020 18300 11026 18312
rect 11517 18309 11529 18312
rect 11563 18309 11575 18343
rect 11517 18303 11575 18309
rect 18417 18343 18475 18349
rect 18417 18309 18429 18343
rect 18463 18340 18475 18343
rect 19426 18340 19432 18352
rect 18463 18312 19432 18340
rect 18463 18309 18475 18312
rect 18417 18303 18475 18309
rect 19426 18300 19432 18312
rect 19484 18340 19490 18352
rect 19484 18312 19656 18340
rect 19484 18300 19490 18312
rect 2038 18232 2044 18284
rect 2096 18272 2102 18284
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 2096 18244 2237 18272
rect 2096 18232 2102 18244
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4120 18244 4292 18272
rect 4120 18232 4126 18244
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18136 2007 18139
rect 2501 18139 2559 18145
rect 2501 18136 2513 18139
rect 1995 18108 2513 18136
rect 1995 18105 2007 18108
rect 1949 18099 2007 18105
rect 2501 18105 2513 18108
rect 2547 18136 2559 18139
rect 2590 18136 2596 18148
rect 2547 18108 2596 18136
rect 2547 18105 2559 18108
rect 2501 18099 2559 18105
rect 2590 18096 2596 18108
rect 2648 18096 2654 18148
rect 2958 18096 2964 18148
rect 3016 18096 3022 18148
rect 4264 18145 4292 18244
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 6089 18275 6147 18281
rect 6089 18272 6101 18275
rect 5408 18244 6101 18272
rect 5408 18232 5414 18244
rect 6089 18241 6101 18244
rect 6135 18241 6147 18275
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 6089 18235 6147 18241
rect 7024 18244 7573 18272
rect 7024 18213 7052 18244
rect 7561 18241 7573 18244
rect 7607 18272 7619 18275
rect 8754 18272 8760 18284
rect 7607 18244 8760 18272
rect 7607 18241 7619 18244
rect 7561 18235 7619 18241
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9631 18244 10272 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18173 7067 18207
rect 7834 18204 7840 18216
rect 7747 18176 7840 18204
rect 7009 18167 7067 18173
rect 7834 18164 7840 18176
rect 7892 18204 7898 18216
rect 9858 18204 9864 18216
rect 7892 18176 8340 18204
rect 9819 18176 9864 18204
rect 7892 18164 7898 18176
rect 4249 18139 4307 18145
rect 4249 18105 4261 18139
rect 4295 18136 4307 18139
rect 4525 18139 4583 18145
rect 4525 18136 4537 18139
rect 4295 18108 4537 18136
rect 4295 18105 4307 18108
rect 4249 18099 4307 18105
rect 4525 18105 4537 18108
rect 4571 18105 4583 18139
rect 4525 18099 4583 18105
rect 8312 18080 8340 18176
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10042 18204 10048 18216
rect 10003 18176 10048 18204
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10244 18204 10272 18244
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 14148 18244 14473 18272
rect 14148 18232 14154 18244
rect 14461 18241 14473 18244
rect 14507 18272 14519 18275
rect 15102 18272 15108 18284
rect 14507 18244 15108 18272
rect 14507 18241 14519 18244
rect 14461 18235 14519 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16485 18275 16543 18281
rect 16485 18272 16497 18275
rect 15988 18244 16497 18272
rect 15988 18232 15994 18244
rect 16485 18241 16497 18244
rect 16531 18272 16543 18275
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 16531 18244 16773 18272
rect 16531 18241 16543 18244
rect 16485 18235 16543 18241
rect 16761 18241 16773 18244
rect 16807 18241 16819 18275
rect 16761 18235 16819 18241
rect 10502 18204 10508 18216
rect 10244 18176 10508 18204
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 19628 18213 19656 18312
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18173 10655 18207
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 10597 18167 10655 18173
rect 16684 18176 18245 18204
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18136 8907 18139
rect 10060 18136 10088 18164
rect 8895 18108 10088 18136
rect 8895 18105 8907 18108
rect 8849 18099 8907 18105
rect 10318 18096 10324 18148
rect 10376 18136 10382 18148
rect 10612 18136 10640 18167
rect 10376 18108 10640 18136
rect 14185 18139 14243 18145
rect 10376 18096 10382 18108
rect 14185 18105 14197 18139
rect 14231 18136 14243 18139
rect 14734 18136 14740 18148
rect 14231 18108 14740 18136
rect 14231 18105 14243 18108
rect 14185 18099 14243 18105
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 15746 18096 15752 18148
rect 15804 18096 15810 18148
rect 8018 18068 8024 18080
rect 7979 18040 8024 18068
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 8294 18068 8300 18080
rect 8255 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 16684 18068 16712 18176
rect 18233 18173 18245 18176
rect 18279 18204 18291 18207
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 18279 18176 18705 18204
rect 18279 18173 18291 18176
rect 18233 18167 18291 18173
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 19613 18207 19671 18213
rect 19613 18173 19625 18207
rect 19659 18173 19671 18207
rect 20438 18204 20444 18216
rect 20399 18176 20444 18204
rect 19613 18167 19671 18173
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 22278 18204 22284 18216
rect 22239 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18204 22342 18216
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22336 18176 22753 18204
rect 22336 18164 22342 18176
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 22741 18167 22799 18173
rect 19058 18068 19064 18080
rect 13136 18040 16712 18068
rect 19019 18040 19064 18068
rect 13136 18028 13142 18040
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 22462 18068 22468 18080
rect 22423 18040 22468 18068
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 1104 17978 24656 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 24656 17978
rect 1104 17904 24656 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2958 17864 2964 17876
rect 2363 17836 2964 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2958 17824 2964 17836
rect 3016 17864 3022 17876
rect 4433 17867 4491 17873
rect 4433 17864 4445 17867
rect 3016 17836 4445 17864
rect 3016 17824 3022 17836
rect 4433 17833 4445 17836
rect 4479 17833 4491 17867
rect 4433 17827 4491 17833
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 8294 17864 8300 17876
rect 8067 17836 8300 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8294 17824 8300 17836
rect 8352 17864 8358 17876
rect 8665 17867 8723 17873
rect 8665 17864 8677 17867
rect 8352 17836 8677 17864
rect 8352 17824 8358 17836
rect 8665 17833 8677 17836
rect 8711 17833 8723 17867
rect 8665 17827 8723 17833
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 10042 17864 10048 17876
rect 9355 17836 10048 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 12066 17864 12072 17876
rect 10827 17836 12072 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 14553 17867 14611 17873
rect 14553 17833 14565 17867
rect 14599 17864 14611 17867
rect 15746 17864 15752 17876
rect 14599 17836 15752 17864
rect 14599 17833 14611 17836
rect 14553 17827 14611 17833
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 18969 17867 19027 17873
rect 18969 17833 18981 17867
rect 19015 17864 19027 17867
rect 19150 17864 19156 17876
rect 19015 17836 19156 17864
rect 19015 17833 19027 17836
rect 18969 17827 19027 17833
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19484 17836 19625 17864
rect 19484 17824 19490 17836
rect 19613 17833 19625 17836
rect 19659 17864 19671 17867
rect 20441 17867 20499 17873
rect 20441 17864 20453 17867
rect 19659 17836 20453 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 20441 17833 20453 17836
rect 20487 17864 20499 17867
rect 20898 17864 20904 17876
rect 20487 17836 20904 17864
rect 20487 17833 20499 17836
rect 20441 17827 20499 17833
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 2096 17768 2605 17796
rect 2096 17756 2102 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 3050 17796 3056 17808
rect 3011 17768 3056 17796
rect 2593 17759 2651 17765
rect 2608 17728 2636 17759
rect 3050 17756 3056 17768
rect 3108 17756 3114 17808
rect 13078 17796 13084 17808
rect 13039 17768 13084 17796
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 13909 17799 13967 17805
rect 13909 17765 13921 17799
rect 13955 17796 13967 17799
rect 14918 17796 14924 17808
rect 13955 17768 14924 17796
rect 13955 17765 13967 17768
rect 13909 17759 13967 17765
rect 14918 17756 14924 17768
rect 14976 17796 14982 17808
rect 14976 17768 16528 17796
rect 14976 17756 14982 17768
rect 16500 17740 16528 17768
rect 22462 17756 22468 17808
rect 22520 17756 22526 17808
rect 3234 17728 3240 17740
rect 2608 17700 3240 17728
rect 3234 17688 3240 17700
rect 3292 17728 3298 17740
rect 3329 17731 3387 17737
rect 3329 17728 3341 17731
rect 3292 17700 3341 17728
rect 3292 17688 3298 17700
rect 3329 17697 3341 17700
rect 3375 17697 3387 17731
rect 3329 17691 3387 17697
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 4614 17728 4620 17740
rect 4295 17700 4620 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 5920 17700 6377 17728
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 5350 17660 5356 17672
rect 4847 17632 5356 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 5920 17592 5948 17700
rect 6365 17697 6377 17700
rect 6411 17728 6423 17731
rect 6822 17728 6828 17740
rect 6411 17700 6828 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 6972 17700 7113 17728
rect 6972 17688 6978 17700
rect 7101 17697 7113 17700
rect 7147 17728 7159 17731
rect 8202 17728 8208 17740
rect 7147 17700 8208 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8570 17728 8576 17740
rect 8527 17700 8576 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9088 17700 9873 17728
rect 9088 17688 9094 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 11480 17700 11529 17728
rect 11480 17688 11486 17700
rect 11517 17697 11529 17700
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 11756 17700 12633 17728
rect 11756 17688 11762 17700
rect 12621 17697 12633 17700
rect 12667 17728 12679 17731
rect 13262 17728 13268 17740
rect 12667 17700 13268 17728
rect 12667 17697 12679 17700
rect 12621 17691 12679 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17697 16175 17731
rect 16482 17728 16488 17740
rect 16443 17700 16488 17728
rect 16117 17691 16175 17697
rect 7466 17660 7472 17672
rect 7427 17632 7472 17660
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12124 17632 12541 17660
rect 12124 17620 12130 17632
rect 12529 17629 12541 17632
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 15473 17663 15531 17669
rect 15473 17660 15485 17663
rect 14056 17632 15485 17660
rect 14056 17620 14062 17632
rect 15473 17629 15485 17632
rect 15519 17629 15531 17663
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15473 17623 15531 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 5368 17564 5948 17592
rect 16132 17592 16160 17691
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 17310 17688 17316 17740
rect 17368 17728 17374 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17368 17700 17693 17728
rect 17368 17688 17374 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 18785 17731 18843 17737
rect 18785 17728 18797 17731
rect 17828 17700 18797 17728
rect 17828 17688 17834 17700
rect 18785 17697 18797 17700
rect 18831 17728 18843 17731
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18831 17700 19257 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 16390 17660 16396 17672
rect 16351 17632 16396 17660
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17660 18291 17663
rect 18966 17660 18972 17672
rect 18279 17632 18972 17660
rect 18279 17629 18291 17632
rect 18233 17623 18291 17629
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 21726 17660 21732 17672
rect 21687 17632 21732 17660
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 22428 17632 23489 17660
rect 22428 17620 22434 17632
rect 23477 17629 23489 17632
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 16132 17564 17080 17592
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5368 17533 5396 17564
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 5040 17496 5365 17524
rect 5040 17484 5046 17496
rect 5353 17493 5365 17496
rect 5399 17493 5411 17527
rect 5353 17487 5411 17493
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9858 17524 9864 17536
rect 9364 17496 9864 17524
rect 9364 17484 9370 17496
rect 9858 17484 9864 17496
rect 9916 17524 9922 17536
rect 10045 17527 10103 17533
rect 10045 17524 10057 17527
rect 9916 17496 10057 17524
rect 9916 17484 9922 17496
rect 10045 17493 10057 17496
rect 10091 17524 10103 17527
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10091 17496 10333 17524
rect 10091 17493 10103 17496
rect 10045 17487 10103 17493
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 11054 17524 11060 17536
rect 11015 17496 11060 17524
rect 10321 17487 10379 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 17052 17533 17080 17564
rect 11701 17527 11759 17533
rect 11701 17524 11713 17527
rect 11572 17496 11713 17524
rect 11572 17484 11578 17496
rect 11701 17493 11713 17496
rect 11747 17493 11759 17527
rect 11701 17487 11759 17493
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 17083 17496 17417 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17405 17493 17417 17496
rect 17451 17524 17463 17527
rect 17494 17524 17500 17536
rect 17451 17496 17500 17524
rect 17451 17493 17463 17496
rect 17405 17487 17463 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17862 17524 17868 17536
rect 17823 17496 17868 17524
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 21048 17496 21097 17524
rect 21048 17484 21054 17496
rect 21085 17493 21097 17496
rect 21131 17524 21143 17527
rect 21818 17524 21824 17536
rect 21131 17496 21824 17524
rect 21131 17493 21143 17496
rect 21085 17487 21143 17493
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 1104 17434 24656 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 24656 17434
rect 1104 17360 24656 17382
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 6089 17323 6147 17329
rect 6089 17320 6101 17323
rect 5500 17292 6101 17320
rect 5500 17280 5506 17292
rect 6089 17289 6101 17292
rect 6135 17320 6147 17323
rect 6914 17320 6920 17332
rect 6135 17292 6920 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 15565 17323 15623 17329
rect 15565 17289 15577 17323
rect 15611 17320 15623 17323
rect 15930 17320 15936 17332
rect 15611 17292 15936 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 16482 17320 16488 17332
rect 16443 17292 16488 17320
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 17310 17320 17316 17332
rect 17271 17292 17316 17320
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 22557 17323 22615 17329
rect 22557 17320 22569 17323
rect 22520 17292 22569 17320
rect 22520 17280 22526 17292
rect 22557 17289 22569 17292
rect 22603 17289 22615 17323
rect 22557 17283 22615 17289
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 14458 17252 14464 17264
rect 13035 17224 14464 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 14458 17212 14464 17224
rect 14516 17212 14522 17264
rect 14734 17212 14740 17264
rect 14792 17252 14798 17264
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 14792 17224 14933 17252
rect 14792 17212 14798 17224
rect 14921 17221 14933 17224
rect 14967 17221 14979 17255
rect 14921 17215 14979 17221
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 21726 17252 21732 17264
rect 20671 17224 21732 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 21726 17212 21732 17224
rect 21784 17252 21790 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21784 17224 22017 17252
rect 21784 17212 21790 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 2406 17184 2412 17196
rect 1903 17156 2412 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 17681 17187 17739 17193
rect 12952 17156 14136 17184
rect 12952 17144 12958 17156
rect 14108 17128 14136 17156
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 18509 17187 18567 17193
rect 18509 17184 18521 17187
rect 17727 17156 18521 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 18509 17153 18521 17156
rect 18555 17184 18567 17187
rect 18598 17184 18604 17196
rect 18555 17156 18604 17184
rect 18555 17153 18567 17156
rect 18509 17147 18567 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 20898 17184 20904 17196
rect 20859 17156 20904 17184
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2133 17119 2191 17125
rect 2133 17116 2145 17119
rect 2096 17088 2145 17116
rect 2096 17076 2102 17088
rect 2133 17085 2145 17088
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4120 17088 4997 17116
rect 4120 17076 4126 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 5350 17116 5356 17128
rect 5311 17088 5356 17116
rect 4985 17079 5043 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6457 17119 6515 17125
rect 6457 17085 6469 17119
rect 6503 17116 6515 17119
rect 6638 17116 6644 17128
rect 6503 17088 6644 17116
rect 6503 17085 6515 17088
rect 6457 17079 6515 17085
rect 6638 17076 6644 17088
rect 6696 17116 6702 17128
rect 7101 17119 7159 17125
rect 7101 17116 7113 17119
rect 6696 17088 7113 17116
rect 6696 17076 6702 17088
rect 7101 17085 7113 17088
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 9364 17088 9413 17116
rect 9364 17076 9370 17088
rect 9401 17085 9413 17088
rect 9447 17085 9459 17119
rect 10042 17116 10048 17128
rect 10003 17088 10048 17116
rect 9401 17079 9459 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 13170 17116 13176 17128
rect 12851 17088 13176 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 13998 17116 14004 17128
rect 13959 17088 14004 17116
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14461 17119 14519 17125
rect 14148 17088 14193 17116
rect 14148 17076 14154 17088
rect 14461 17085 14473 17119
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17116 14611 17119
rect 14918 17116 14924 17128
rect 14599 17088 14924 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 3142 17008 3148 17060
rect 3200 17008 3206 17060
rect 3694 17008 3700 17060
rect 3752 17048 3758 17060
rect 4157 17051 4215 17057
rect 4157 17048 4169 17051
rect 3752 17020 4169 17048
rect 3752 17008 3758 17020
rect 4157 17017 4169 17020
rect 4203 17048 4215 17051
rect 5368 17048 5396 17076
rect 4203 17020 5396 17048
rect 4203 17017 4215 17020
rect 4157 17011 4215 17017
rect 6086 17008 6092 17060
rect 6144 17048 6150 17060
rect 7009 17051 7067 17057
rect 7009 17048 7021 17051
rect 6144 17020 7021 17048
rect 6144 17008 6150 17020
rect 7009 17017 7021 17020
rect 7055 17017 7067 17051
rect 7009 17011 7067 17017
rect 10778 17008 10784 17060
rect 10836 17008 10842 17060
rect 14476 17048 14504 17079
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17116 16727 17119
rect 17494 17116 17500 17128
rect 16715 17088 17500 17116
rect 16715 17085 16727 17088
rect 16669 17079 16727 17085
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 18230 17116 18236 17128
rect 18191 17088 18236 17116
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 21082 17116 21088 17128
rect 21043 17088 21088 17116
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 21174 17076 21180 17128
rect 21232 17116 21238 17128
rect 21545 17119 21603 17125
rect 21545 17116 21557 17119
rect 21232 17088 21557 17116
rect 21232 17076 21238 17088
rect 21545 17085 21557 17088
rect 21591 17085 21603 17119
rect 21545 17079 21603 17085
rect 21637 17119 21695 17125
rect 21637 17085 21649 17119
rect 21683 17116 21695 17119
rect 22646 17116 22652 17128
rect 21683 17088 22652 17116
rect 21683 17085 21695 17088
rect 21637 17079 21695 17085
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 14826 17048 14832 17060
rect 14476 17020 14832 17048
rect 14826 17008 14832 17020
rect 14884 17048 14890 17060
rect 16390 17048 16396 17060
rect 14884 17020 16396 17048
rect 14884 17008 14890 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 18966 17008 18972 17060
rect 19024 17008 19030 17060
rect 20254 17048 20260 17060
rect 20215 17020 20260 17048
rect 20254 17008 20260 17020
rect 20312 17008 20318 17060
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4614 16980 4620 16992
rect 4571 16952 4620 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4614 16940 4620 16952
rect 4672 16980 4678 16992
rect 5074 16980 5080 16992
rect 4672 16952 5080 16980
rect 4672 16940 4678 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 8570 16980 8576 16992
rect 8531 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 11422 16980 11428 16992
rect 10284 16952 11428 16980
rect 10284 16940 10290 16952
rect 11422 16940 11428 16952
rect 11480 16980 11486 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 11480 16952 11529 16980
rect 11480 16940 11486 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 12066 16980 12072 16992
rect 12027 16952 12072 16980
rect 11517 16943 11575 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 21450 16940 21456 16992
rect 21508 16980 21514 16992
rect 22922 16980 22928 16992
rect 21508 16952 22928 16980
rect 21508 16940 21514 16952
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 1104 16890 24656 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 24656 16890
rect 1104 16816 24656 16838
rect 2225 16779 2283 16785
rect 2225 16745 2237 16779
rect 2271 16776 2283 16779
rect 3142 16776 3148 16788
rect 2271 16748 3148 16776
rect 2271 16745 2283 16748
rect 2225 16739 2283 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3234 16736 3240 16788
rect 3292 16776 3298 16788
rect 3694 16776 3700 16788
rect 3292 16748 3337 16776
rect 3655 16748 3700 16776
rect 3292 16736 3298 16748
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 6822 16776 6828 16788
rect 6783 16748 6828 16776
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7285 16779 7343 16785
rect 7285 16745 7297 16779
rect 7331 16776 7343 16779
rect 8018 16776 8024 16788
rect 7331 16748 8024 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9306 16776 9312 16788
rect 9267 16748 9312 16776
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 13541 16779 13599 16785
rect 13541 16745 13553 16779
rect 13587 16776 13599 16779
rect 13998 16776 14004 16788
rect 13587 16748 14004 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 14148 16748 14197 16776
rect 14148 16736 14154 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14826 16776 14832 16788
rect 14787 16748 14832 16776
rect 14185 16739 14243 16745
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 15488 16748 17877 16776
rect 1670 16668 1676 16720
rect 1728 16708 1734 16720
rect 2314 16708 2320 16720
rect 1728 16680 2320 16708
rect 1728 16668 1734 16680
rect 2314 16668 2320 16680
rect 2372 16708 2378 16720
rect 2869 16711 2927 16717
rect 2869 16708 2881 16711
rect 2372 16680 2881 16708
rect 2372 16668 2378 16680
rect 2869 16677 2881 16680
rect 2915 16677 2927 16711
rect 2869 16671 2927 16677
rect 4801 16711 4859 16717
rect 4801 16677 4813 16711
rect 4847 16708 4859 16711
rect 4847 16680 6132 16708
rect 4847 16677 4859 16680
rect 4801 16671 4859 16677
rect 6104 16652 6132 16680
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 11057 16711 11115 16717
rect 11057 16708 11069 16711
rect 10836 16680 11069 16708
rect 10836 16668 10842 16680
rect 11057 16677 11069 16680
rect 11103 16677 11115 16711
rect 11057 16671 11115 16677
rect 11514 16668 11520 16720
rect 11572 16668 11578 16720
rect 13909 16711 13967 16717
rect 13909 16677 13921 16711
rect 13955 16708 13967 16711
rect 14844 16708 14872 16736
rect 13955 16680 14872 16708
rect 13955 16677 13967 16680
rect 13909 16671 13967 16677
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5353 16643 5411 16649
rect 5353 16640 5365 16643
rect 5040 16612 5365 16640
rect 5040 16600 5046 16612
rect 5353 16609 5365 16612
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 5902 16640 5908 16652
rect 5500 16612 5545 16640
rect 5863 16612 5908 16640
rect 5500 16600 5506 16612
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 6086 16640 6092 16652
rect 6047 16612 6092 16640
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 8570 16640 8576 16652
rect 8483 16612 8576 16640
rect 8570 16600 8576 16612
rect 8628 16640 8634 16652
rect 9858 16640 9864 16652
rect 8628 16612 9864 16640
rect 8628 16600 8634 16612
rect 9858 16600 9864 16612
rect 9916 16640 9922 16652
rect 9916 16612 10364 16640
rect 9916 16600 9922 16612
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2498 16572 2504 16584
rect 1719 16544 2504 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 4890 16464 4896 16516
rect 4948 16504 4954 16516
rect 6273 16507 6331 16513
rect 6273 16504 6285 16507
rect 4948 16476 6285 16504
rect 4948 16464 4954 16476
rect 6273 16473 6285 16476
rect 6319 16473 6331 16507
rect 6273 16467 6331 16473
rect 1670 16396 1676 16448
rect 1728 16436 1734 16448
rect 2501 16439 2559 16445
rect 2501 16436 2513 16439
rect 1728 16408 2513 16436
rect 1728 16396 1734 16408
rect 2501 16405 2513 16408
rect 2547 16405 2559 16439
rect 2501 16399 2559 16405
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 4120 16408 4353 16436
rect 4120 16396 4126 16408
rect 4341 16405 4353 16408
rect 4387 16405 4399 16439
rect 8754 16436 8760 16448
rect 8715 16408 8760 16436
rect 4341 16399 4399 16405
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 10045 16439 10103 16445
rect 10045 16405 10057 16439
rect 10091 16436 10103 16439
rect 10226 16436 10232 16448
rect 10091 16408 10232 16436
rect 10091 16405 10103 16408
rect 10045 16399 10103 16405
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 10336 16436 10364 16612
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15488 16649 15516 16748
rect 17865 16745 17877 16748
rect 17911 16776 17923 16779
rect 18230 16776 18236 16788
rect 17911 16748 18236 16776
rect 17911 16745 17923 16748
rect 17865 16739 17923 16745
rect 18230 16736 18236 16748
rect 18288 16776 18294 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18288 16748 18613 16776
rect 18288 16736 18294 16748
rect 18601 16745 18613 16748
rect 18647 16745 18659 16779
rect 18601 16739 18659 16745
rect 18966 16736 18972 16788
rect 19024 16776 19030 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 19024 16748 19257 16776
rect 19024 16736 19030 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 19245 16739 19303 16745
rect 16482 16668 16488 16720
rect 16540 16668 16546 16720
rect 17494 16708 17500 16720
rect 17455 16680 17500 16708
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 20165 16711 20223 16717
rect 20165 16677 20177 16711
rect 20211 16708 20223 16711
rect 20438 16708 20444 16720
rect 20211 16680 20444 16708
rect 20211 16677 20223 16680
rect 20165 16671 20223 16677
rect 20438 16668 20444 16680
rect 20496 16708 20502 16720
rect 21082 16708 21088 16720
rect 20496 16680 21088 16708
rect 20496 16668 20502 16680
rect 21082 16668 21088 16680
rect 21140 16708 21146 16720
rect 21637 16711 21695 16717
rect 21637 16708 21649 16711
rect 21140 16680 21649 16708
rect 21140 16668 21146 16680
rect 21637 16677 21649 16680
rect 21683 16677 21695 16711
rect 21637 16671 21695 16677
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15160 16612 15485 16640
rect 15160 16600 15166 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 19058 16640 19064 16652
rect 18971 16612 19064 16640
rect 15473 16603 15531 16609
rect 19058 16600 19064 16612
rect 19116 16640 19122 16652
rect 19426 16640 19432 16652
rect 19116 16612 19432 16640
rect 19116 16600 19122 16612
rect 19426 16600 19432 16612
rect 19484 16600 19490 16652
rect 22278 16640 22284 16652
rect 22239 16612 22284 16640
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22646 16640 22652 16652
rect 22607 16612 22652 16640
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16572 10839 16575
rect 11054 16572 11060 16584
rect 10827 16544 11060 16572
rect 10827 16541 10839 16544
rect 10781 16535 10839 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 12802 16572 12808 16584
rect 12763 16544 12808 16572
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 22370 16572 22376 16584
rect 22331 16544 22376 16572
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 22554 16572 22560 16584
rect 22515 16544 22560 16572
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 18325 16507 18383 16513
rect 18325 16473 18337 16507
rect 18371 16504 18383 16507
rect 18782 16504 18788 16516
rect 18371 16476 18788 16504
rect 18371 16473 18383 16476
rect 18325 16467 18383 16473
rect 18782 16464 18788 16476
rect 18840 16464 18846 16516
rect 13170 16436 13176 16448
rect 10336 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 20530 16436 20536 16448
rect 20491 16408 20536 16436
rect 20530 16396 20536 16408
rect 20588 16396 20594 16448
rect 21174 16436 21180 16448
rect 21135 16408 21180 16436
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 1104 16346 24656 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 24656 16346
rect 1104 16272 24656 16294
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6144 16204 6193 16232
rect 6144 16192 6150 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 9858 16232 9864 16244
rect 9819 16204 9864 16232
rect 6181 16195 6239 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10229 16235 10287 16241
rect 10229 16201 10241 16235
rect 10275 16232 10287 16235
rect 11514 16232 11520 16244
rect 10275 16204 11520 16232
rect 10275 16201 10287 16204
rect 10229 16195 10287 16201
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 12805 16235 12863 16241
rect 12805 16201 12817 16235
rect 12851 16232 12863 16235
rect 12894 16232 12900 16244
rect 12851 16204 12900 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 15102 16232 15108 16244
rect 15063 16204 15108 16232
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15841 16235 15899 16241
rect 15841 16201 15853 16235
rect 15887 16232 15899 16235
rect 16482 16232 16488 16244
rect 15887 16204 16488 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 16577 16235 16635 16241
rect 16577 16201 16589 16235
rect 16623 16232 16635 16235
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 16623 16204 16865 16232
rect 16623 16201 16635 16204
rect 16577 16195 16635 16201
rect 16853 16201 16865 16204
rect 16899 16232 16911 16235
rect 17770 16232 17776 16244
rect 16899 16204 17776 16232
rect 16899 16201 16911 16204
rect 16853 16195 16911 16201
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 20530 16192 20536 16244
rect 20588 16232 20594 16244
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 20588 16204 21005 16232
rect 20588 16192 20594 16204
rect 20993 16201 21005 16204
rect 21039 16232 21051 16235
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 21039 16204 22477 16232
rect 21039 16201 21051 16204
rect 20993 16195 21051 16201
rect 22465 16201 22477 16204
rect 22511 16232 22523 16235
rect 22646 16232 22652 16244
rect 22511 16204 22652 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 21361 16167 21419 16173
rect 21361 16164 21373 16167
rect 21232 16136 21373 16164
rect 21232 16124 21238 16136
rect 21361 16133 21373 16136
rect 21407 16164 21419 16167
rect 22554 16164 22560 16176
rect 21407 16136 22560 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 4062 16096 4068 16108
rect 3975 16068 4068 16096
rect 4062 16056 4068 16068
rect 4120 16096 4126 16108
rect 5902 16096 5908 16108
rect 4120 16068 5908 16096
rect 4120 16056 4126 16068
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 16028 4491 16031
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4479 16000 5181 16028
rect 4479 15997 4491 16000
rect 4433 15991 4491 15997
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5350 16028 5356 16040
rect 5311 16000 5356 16028
rect 5169 15991 5227 15997
rect 2590 15920 2596 15972
rect 2648 15920 2654 15972
rect 5184 15960 5212 15991
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5736 16037 5764 16068
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 7466 16096 7472 16108
rect 7427 16068 7472 16096
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 8478 16056 8484 16108
rect 8536 16096 8542 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 8536 16068 10517 16096
rect 8536 16056 8542 16068
rect 10505 16065 10517 16068
rect 10551 16096 10563 16099
rect 11146 16096 11152 16108
rect 10551 16068 11152 16096
rect 10551 16065 10563 16068
rect 10505 16059 10563 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15746 16096 15752 16108
rect 15519 16068 15752 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15746 16056 15752 16068
rect 15804 16096 15810 16108
rect 19242 16096 19248 16108
rect 15804 16068 19248 16096
rect 15804 16056 15810 16068
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 21729 16099 21787 16105
rect 21729 16065 21741 16099
rect 21775 16096 21787 16099
rect 22370 16096 22376 16108
rect 21775 16068 22376 16096
rect 21775 16065 21787 16068
rect 21729 16059 21787 16065
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 6086 16028 6092 16040
rect 5859 16000 6092 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6086 15988 6092 16000
rect 6144 15988 6150 16040
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 16028 9275 16031
rect 10134 16028 10140 16040
rect 9263 16000 10140 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 11103 16000 12633 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 12621 15997 12633 16000
rect 12667 16028 12679 16031
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 12667 16000 13093 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13081 15997 13093 16000
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 6638 15960 6644 15972
rect 5184 15932 6644 15960
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 8018 15920 8024 15972
rect 8076 15920 8082 15972
rect 10410 15920 10416 15972
rect 10468 15960 10474 15972
rect 10612 15960 10640 15991
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13228 16000 14105 16028
rect 13228 15988 13234 16000
rect 14093 15997 14105 16000
rect 14139 16028 14151 16031
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 14139 16000 14565 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 16577 16031 16635 16037
rect 16577 16028 16589 16031
rect 16347 16000 16589 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16577 15997 16589 16000
rect 16623 15997 16635 16031
rect 18230 16028 18236 16040
rect 18191 16000 18236 16028
rect 16577 15991 16635 15997
rect 11333 15963 11391 15969
rect 11333 15960 11345 15963
rect 10468 15932 11345 15960
rect 10468 15920 10474 15932
rect 11333 15929 11345 15932
rect 11379 15929 11391 15963
rect 16316 15960 16344 15991
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 16028 20683 16031
rect 22278 16028 22284 16040
rect 20671 16000 22284 16028
rect 20671 15997 20683 16000
rect 20625 15991 20683 15997
rect 22278 15988 22284 16000
rect 22336 16028 22342 16040
rect 22649 16031 22707 16037
rect 22649 16028 22661 16031
rect 22336 16000 22661 16028
rect 22336 15988 22342 16000
rect 22649 15997 22661 16000
rect 22695 16028 22707 16031
rect 22695 16000 23152 16028
rect 22695 15997 22707 16000
rect 22649 15991 22707 15997
rect 11333 15923 11391 15929
rect 14292 15932 16344 15960
rect 18509 15963 18567 15969
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 11112 15864 11713 15892
rect 11112 15852 11118 15864
rect 11701 15861 11713 15864
rect 11747 15861 11759 15895
rect 11701 15855 11759 15861
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14292 15901 14320 15932
rect 18509 15929 18521 15963
rect 18555 15960 18567 15963
rect 18782 15960 18788 15972
rect 18555 15932 18788 15960
rect 18555 15929 18567 15932
rect 18509 15923 18567 15929
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 20257 15963 20315 15969
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 14240 15864 14289 15892
rect 14240 15852 14246 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 17681 15895 17739 15901
rect 17681 15861 17693 15895
rect 17727 15892 17739 15895
rect 17862 15892 17868 15904
rect 17727 15864 17868 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 17862 15852 17868 15864
rect 17920 15892 17926 15904
rect 18984 15892 19012 15960
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 20898 15960 20904 15972
rect 20303 15932 20904 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 23124 15901 23152 16000
rect 17920 15864 19012 15892
rect 23109 15895 23167 15901
rect 17920 15852 17926 15864
rect 23109 15861 23121 15895
rect 23155 15892 23167 15895
rect 23382 15892 23388 15904
rect 23155 15864 23388 15892
rect 23155 15861 23167 15864
rect 23109 15855 23167 15861
rect 23382 15852 23388 15864
rect 23440 15852 23446 15904
rect 1104 15802 24656 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 24656 15802
rect 1104 15728 24656 15750
rect 7285 15691 7343 15697
rect 7285 15657 7297 15691
rect 7331 15688 7343 15691
rect 7466 15688 7472 15700
rect 7331 15660 7472 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8570 15688 8576 15700
rect 8531 15660 8576 15688
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 11146 15648 11152 15660
rect 11204 15688 11210 15700
rect 12526 15688 12532 15700
rect 11204 15660 12532 15688
rect 11204 15648 11210 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 18601 15691 18659 15697
rect 18601 15657 18613 15691
rect 18647 15688 18659 15691
rect 20990 15688 20996 15700
rect 18647 15660 20996 15688
rect 18647 15657 18659 15660
rect 18601 15651 18659 15657
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 2590 15620 2596 15632
rect 2332 15592 2596 15620
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 1854 15552 1860 15564
rect 1811 15524 1860 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 1854 15512 1860 15524
rect 1912 15552 1918 15564
rect 2222 15552 2228 15564
rect 1912 15524 2228 15552
rect 1912 15512 1918 15524
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 2332 15561 2360 15592
rect 2590 15580 2596 15592
rect 2648 15620 2654 15632
rect 3237 15623 3295 15629
rect 3237 15620 3249 15623
rect 2648 15592 3249 15620
rect 2648 15580 2654 15592
rect 3237 15589 3249 15592
rect 3283 15589 3295 15623
rect 4890 15620 4896 15632
rect 4851 15592 4896 15620
rect 3237 15583 3295 15589
rect 4890 15580 4896 15592
rect 4948 15580 4954 15632
rect 5534 15580 5540 15632
rect 5592 15580 5598 15632
rect 6638 15620 6644 15632
rect 6599 15592 6644 15620
rect 6638 15580 6644 15592
rect 6696 15580 6702 15632
rect 16945 15623 17003 15629
rect 16945 15589 16957 15623
rect 16991 15620 17003 15623
rect 17034 15620 17040 15632
rect 16991 15592 17040 15620
rect 16991 15589 17003 15592
rect 16945 15583 17003 15589
rect 17034 15580 17040 15592
rect 17092 15620 17098 15632
rect 20254 15620 20260 15632
rect 17092 15592 20260 15620
rect 17092 15580 17098 15592
rect 20254 15580 20260 15592
rect 20312 15580 20318 15632
rect 22554 15620 22560 15632
rect 22515 15592 22560 15620
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15521 2375 15555
rect 2498 15552 2504 15564
rect 2459 15524 2504 15552
rect 2317 15515 2375 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 10226 15552 10232 15564
rect 10187 15524 10232 15552
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 13078 15552 13084 15564
rect 13039 15524 13084 15552
rect 13078 15512 13084 15524
rect 13136 15512 13142 15564
rect 15930 15552 15936 15564
rect 15891 15524 15936 15552
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 20622 15552 20628 15564
rect 19567 15524 20628 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15552 21327 15555
rect 21910 15552 21916 15564
rect 21315 15524 21916 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 22370 15512 22376 15564
rect 22428 15552 22434 15564
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 22428 15524 22661 15552
rect 22428 15512 22434 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 6270 15484 6276 15496
rect 4663 15456 6276 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 6270 15444 6276 15456
rect 6328 15484 6334 15496
rect 7006 15484 7012 15496
rect 6328 15456 7012 15484
rect 6328 15444 6334 15456
rect 7006 15444 7012 15456
rect 7064 15484 7070 15496
rect 7190 15484 7196 15496
rect 7064 15456 7196 15484
rect 7064 15444 7070 15456
rect 7190 15444 7196 15456
rect 7248 15484 7254 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7248 15456 7573 15484
rect 7248 15444 7254 15456
rect 7561 15453 7573 15456
rect 7607 15453 7619 15487
rect 15838 15484 15844 15496
rect 15799 15456 15844 15484
rect 7561 15447 7619 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 2685 15419 2743 15425
rect 2685 15416 2697 15419
rect 2556 15388 2697 15416
rect 2556 15376 2562 15388
rect 2685 15385 2697 15388
rect 2731 15385 2743 15419
rect 2685 15379 2743 15385
rect 14826 15376 14832 15428
rect 14884 15416 14890 15428
rect 19444 15416 19472 15447
rect 20257 15419 20315 15425
rect 20257 15416 20269 15419
rect 14884 15388 20269 15416
rect 14884 15376 14890 15388
rect 20257 15385 20269 15388
rect 20303 15416 20315 15419
rect 21192 15416 21220 15447
rect 22005 15419 22063 15425
rect 22005 15416 22017 15419
rect 20303 15388 22017 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 22005 15385 22017 15388
rect 22051 15385 22063 15419
rect 22005 15379 22063 15385
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 3605 15351 3663 15357
rect 3605 15348 3617 15351
rect 1728 15320 3617 15348
rect 1728 15308 1734 15320
rect 3605 15317 3617 15320
rect 3651 15317 3663 15351
rect 3605 15311 3663 15317
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 5442 15348 5448 15360
rect 4387 15320 5448 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 10413 15351 10471 15357
rect 10413 15317 10425 15351
rect 10459 15348 10471 15351
rect 10594 15348 10600 15360
rect 10459 15320 10600 15348
rect 10459 15317 10471 15320
rect 10413 15311 10471 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 12575 15320 13185 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13173 15317 13185 15320
rect 13219 15348 13231 15351
rect 13538 15348 13544 15360
rect 13219 15320 13544 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 18141 15351 18199 15357
rect 18141 15317 18153 15351
rect 18187 15348 18199 15351
rect 18506 15348 18512 15360
rect 18187 15320 18512 15348
rect 18187 15317 18199 15320
rect 18141 15311 18199 15317
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 19153 15351 19211 15357
rect 19153 15317 19165 15351
rect 19199 15348 19211 15351
rect 19426 15348 19432 15360
rect 19199 15320 19432 15348
rect 19199 15317 19211 15320
rect 19153 15311 19211 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19705 15351 19763 15357
rect 19705 15317 19717 15351
rect 19751 15348 19763 15351
rect 19886 15348 19892 15360
rect 19751 15320 19892 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 1104 15258 24656 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 24656 15258
rect 1104 15184 24656 15206
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4890 15144 4896 15156
rect 4755 15116 4896 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 10226 15144 10232 15156
rect 10187 15116 10232 15144
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 15565 15147 15623 15153
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 15838 15144 15844 15156
rect 15611 15116 15844 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 15838 15104 15844 15116
rect 15896 15104 15902 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 18414 15144 18420 15156
rect 17727 15116 18420 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 22833 15147 22891 15153
rect 22833 15144 22845 15147
rect 22428 15116 22845 15144
rect 22428 15104 22434 15116
rect 22833 15113 22845 15116
rect 22879 15113 22891 15147
rect 22833 15107 22891 15113
rect 3602 15036 3608 15088
rect 3660 15076 3666 15088
rect 5261 15079 5319 15085
rect 5261 15076 5273 15079
rect 3660 15048 5273 15076
rect 3660 15036 3666 15048
rect 5261 15045 5273 15048
rect 5307 15045 5319 15079
rect 5261 15039 5319 15045
rect 11701 15079 11759 15085
rect 11701 15045 11713 15079
rect 11747 15076 11759 15079
rect 18432 15076 18460 15104
rect 11747 15048 13400 15076
rect 18432 15048 22416 15076
rect 11747 15045 11759 15048
rect 11701 15039 11759 15045
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2498 15008 2504 15020
rect 1995 14980 2504 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 9030 15008 9036 15020
rect 8991 14980 9036 15008
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 13078 15008 13084 15020
rect 12115 14980 13084 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13372 14952 13400 15048
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 13648 14980 14473 15008
rect 2038 14900 2044 14952
rect 2096 14940 2102 14952
rect 2225 14943 2283 14949
rect 2225 14940 2237 14943
rect 2096 14912 2237 14940
rect 2096 14900 2102 14912
rect 2225 14909 2237 14912
rect 2271 14909 2283 14943
rect 2225 14903 2283 14909
rect 3602 14900 3608 14952
rect 3660 14900 3666 14952
rect 5074 14940 5080 14952
rect 4987 14912 5080 14940
rect 5074 14900 5080 14912
rect 5132 14940 5138 14952
rect 5626 14940 5632 14952
rect 5132 14912 5632 14940
rect 5132 14900 5138 14912
rect 5626 14900 5632 14912
rect 5684 14940 5690 14952
rect 5997 14943 6055 14949
rect 5997 14940 6009 14943
rect 5684 14912 6009 14940
rect 5684 14900 5690 14912
rect 5997 14909 6009 14912
rect 6043 14940 6055 14943
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 6043 14912 7481 14940
rect 6043 14909 6055 14912
rect 5997 14903 6055 14909
rect 7469 14909 7481 14912
rect 7515 14940 7527 14943
rect 7515 14912 8064 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14872 4307 14875
rect 4338 14872 4344 14884
rect 4295 14844 4344 14872
rect 4295 14841 4307 14844
rect 4249 14835 4307 14841
rect 4338 14832 4344 14844
rect 4396 14832 4402 14884
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 7834 14872 7840 14884
rect 7147 14844 7840 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 7650 14804 7656 14816
rect 7611 14776 7656 14804
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 8036 14813 8064 14912
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 8628 14912 9321 14940
rect 8628 14900 8634 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12860 14912 13277 14940
rect 12860 14900 12866 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13280 14872 13308 14903
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 13648 14949 13676 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 22388 14952 22416 15048
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13412 14912 13645 14940
rect 13412 14900 13418 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13633 14903 13691 14909
rect 13786 14912 14197 14940
rect 13786 14872 13814 14912
rect 14185 14909 14197 14912
rect 14231 14940 14243 14943
rect 14550 14940 14556 14952
rect 14231 14912 14556 14940
rect 14231 14909 14243 14912
rect 14185 14903 14243 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 17034 14940 17040 14952
rect 16995 14912 17040 14940
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 18414 14940 18420 14952
rect 18375 14912 18420 14940
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18564 14912 18889 14940
rect 18564 14900 18570 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 20898 14940 20904 14952
rect 20859 14912 20904 14940
rect 18877 14903 18935 14909
rect 20898 14900 20904 14912
rect 20956 14900 20962 14952
rect 22370 14940 22376 14952
rect 22283 14912 22376 14940
rect 22370 14900 22376 14912
rect 22428 14940 22434 14952
rect 23201 14943 23259 14949
rect 23201 14940 23213 14943
rect 22428 14912 23213 14940
rect 22428 14900 22434 14912
rect 23201 14909 23213 14912
rect 23247 14909 23259 14943
rect 23201 14903 23259 14909
rect 16390 14872 16396 14884
rect 13280 14844 13814 14872
rect 16351 14844 16396 14872
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 19242 14832 19248 14884
rect 19300 14832 19306 14884
rect 20254 14832 20260 14884
rect 20312 14872 20318 14884
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 20312 14844 20821 14872
rect 20312 14832 20318 14844
rect 20809 14841 20821 14844
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8754 14804 8760 14816
rect 8067 14776 8760 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8754 14764 8760 14776
rect 8812 14804 8818 14816
rect 10042 14804 10048 14816
rect 8812 14776 10048 14804
rect 8812 14764 8818 14776
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 12710 14804 12716 14816
rect 12671 14776 12716 14804
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 15930 14804 15936 14816
rect 15891 14776 15936 14804
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 22186 14764 22192 14816
rect 22244 14804 22250 14816
rect 22557 14807 22615 14813
rect 22557 14804 22569 14807
rect 22244 14776 22569 14804
rect 22244 14764 22250 14776
rect 22557 14773 22569 14776
rect 22603 14773 22615 14807
rect 22557 14767 22615 14773
rect 1104 14714 24656 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 24656 14714
rect 1104 14640 24656 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3602 14600 3608 14612
rect 3191 14572 3608 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 5626 14600 5632 14612
rect 5587 14572 5632 14600
rect 5626 14560 5632 14572
rect 5684 14560 5690 14612
rect 8478 14600 8484 14612
rect 8439 14572 8484 14600
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 13228 14572 13369 14600
rect 13228 14560 13234 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13357 14563 13415 14569
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14458 14600 14464 14612
rect 14415 14572 14464 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14458 14560 14464 14572
rect 14516 14600 14522 14612
rect 14516 14572 16252 14600
rect 14516 14560 14522 14572
rect 4065 14535 4123 14541
rect 2332 14504 2728 14532
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14433 2283 14467
rect 2225 14427 2283 14433
rect 2240 14328 2268 14427
rect 2332 14405 2360 14504
rect 2590 14464 2596 14476
rect 2551 14436 2596 14464
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 2700 14464 2728 14504
rect 4065 14501 4077 14535
rect 4111 14532 4123 14535
rect 4249 14535 4307 14541
rect 4249 14532 4261 14535
rect 4111 14504 4261 14532
rect 4111 14501 4123 14504
rect 4065 14495 4123 14501
rect 4249 14501 4261 14504
rect 4295 14501 4307 14535
rect 4249 14495 4307 14501
rect 11790 14492 11796 14544
rect 11848 14492 11854 14544
rect 14918 14532 14924 14544
rect 14831 14504 14924 14532
rect 14918 14492 14924 14504
rect 14976 14532 14982 14544
rect 15102 14532 15108 14544
rect 14976 14504 15108 14532
rect 14976 14492 14982 14504
rect 15102 14492 15108 14504
rect 15160 14532 15166 14544
rect 15160 14504 15516 14532
rect 16224 14504 16252 14572
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 18840 14572 19809 14600
rect 18840 14560 18846 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 15160 14492 15166 14504
rect 4338 14464 4344 14476
rect 2700 14436 4344 14464
rect 4338 14424 4344 14436
rect 4396 14464 4402 14476
rect 4893 14467 4951 14473
rect 4893 14464 4905 14467
rect 4396 14436 4905 14464
rect 4396 14424 4402 14436
rect 4893 14433 4905 14436
rect 4939 14464 4951 14467
rect 4982 14464 4988 14476
rect 4939 14436 4988 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7524 14436 7573 14464
rect 7524 14424 7530 14436
rect 7561 14433 7573 14436
rect 7607 14433 7619 14467
rect 7926 14464 7932 14476
rect 7839 14436 7932 14464
rect 7561 14427 7619 14433
rect 7926 14424 7932 14436
rect 7984 14464 7990 14476
rect 9674 14464 9680 14476
rect 7984 14436 9680 14464
rect 7984 14424 7990 14436
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10042 14464 10048 14476
rect 9955 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10686 14464 10692 14476
rect 10100 14436 10692 14464
rect 10100 14424 10106 14436
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 14182 14464 14188 14476
rect 14143 14436 14188 14464
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 15488 14473 15516 14504
rect 19150 14492 19156 14544
rect 19208 14532 19214 14544
rect 19208 14504 19564 14532
rect 19208 14492 19214 14504
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 2406 14396 2412 14408
rect 2363 14368 2412 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2498 14356 2504 14408
rect 2556 14396 2562 14408
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2556 14368 3433 14396
rect 2556 14356 2562 14368
rect 3421 14365 3433 14368
rect 3467 14396 3479 14399
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3467 14368 4077 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7742 14396 7748 14408
rect 7699 14368 7748 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 11054 14396 11060 14408
rect 10967 14368 11060 14396
rect 7837 14359 7895 14365
rect 2774 14328 2780 14340
rect 2240 14300 2780 14328
rect 2774 14288 2780 14300
rect 2832 14288 2838 14340
rect 6641 14331 6699 14337
rect 6641 14297 6653 14331
rect 6687 14328 6699 14331
rect 7852 14328 7880 14359
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11330 14396 11336 14408
rect 11291 14368 11336 14396
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 8018 14328 8024 14340
rect 6687 14300 8024 14328
rect 6687 14297 6699 14300
rect 6641 14291 6699 14297
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10689 14331 10747 14337
rect 10689 14328 10701 14331
rect 9916 14300 10701 14328
rect 9916 14288 9922 14300
rect 10689 14297 10701 14300
rect 10735 14328 10747 14331
rect 11072 14328 11100 14356
rect 10735 14300 11100 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 6270 14260 6276 14272
rect 6231 14232 6276 14260
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 10226 14260 10232 14272
rect 10187 14232 10232 14260
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 15488 14260 15516 14427
rect 18506 14424 18512 14476
rect 18564 14464 18570 14476
rect 18782 14464 18788 14476
rect 18564 14436 18788 14464
rect 18564 14424 18570 14436
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 19334 14464 19340 14476
rect 19295 14436 19340 14464
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 19536 14473 19564 14504
rect 22186 14492 22192 14544
rect 22244 14492 22250 14544
rect 23382 14532 23388 14544
rect 23343 14504 23388 14532
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 20254 14464 20260 14476
rect 19567 14436 20260 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 16114 14356 16120 14408
rect 16172 14396 16178 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 16172 14368 17509 14396
rect 16172 14356 16178 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14396 18199 14399
rect 18414 14396 18420 14408
rect 18187 14368 18420 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 18414 14356 18420 14368
rect 18472 14396 18478 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18472 14368 18613 14396
rect 18472 14356 18478 14368
rect 18601 14365 18613 14368
rect 18647 14396 18659 14399
rect 18874 14396 18880 14408
rect 18647 14368 18880 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 21358 14396 21364 14408
rect 21319 14368 21364 14396
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 22094 14396 22100 14408
rect 21683 14368 22100 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 17218 14260 17224 14272
rect 15488 14232 17224 14260
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20441 14263 20499 14269
rect 20441 14260 20453 14263
rect 20036 14232 20453 14260
rect 20036 14220 20042 14232
rect 20441 14229 20453 14232
rect 20487 14260 20499 14263
rect 20898 14260 20904 14272
rect 20487 14232 20904 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 1104 14170 24656 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 24656 14170
rect 1104 14096 24656 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1765 14059 1823 14065
rect 1765 14056 1777 14059
rect 1728 14028 1777 14056
rect 1728 14016 1734 14028
rect 1765 14025 1777 14028
rect 1811 14025 1823 14059
rect 4982 14056 4988 14068
rect 4943 14028 4988 14056
rect 1765 14019 1823 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 7524 14028 9321 14056
rect 7524 14016 7530 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 4080 13960 5733 13988
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 2682 13920 2688 13932
rect 2096 13892 2688 13920
rect 2096 13880 2102 13892
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 4080 13864 4108 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 6089 13991 6147 13997
rect 6089 13957 6101 13991
rect 6135 13988 6147 13991
rect 6135 13960 7144 13988
rect 6135 13957 6147 13960
rect 6089 13951 6147 13957
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6914 13920 6920 13932
rect 6328 13892 6920 13920
rect 6328 13880 6334 13892
rect 6914 13880 6920 13892
rect 6972 13920 6978 13932
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6972 13892 7021 13920
rect 6972 13880 6978 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7116 13920 7144 13960
rect 7374 13920 7380 13932
rect 7116 13892 7380 13920
rect 7009 13883 7067 13889
rect 7374 13880 7380 13892
rect 7432 13920 7438 13932
rect 7742 13920 7748 13932
rect 7432 13892 7748 13920
rect 7432 13880 7438 13892
rect 7742 13880 7748 13892
rect 7800 13920 7806 13932
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 7800 13892 9045 13920
rect 7800 13880 7806 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13852 1639 13855
rect 2130 13852 2136 13864
rect 1627 13824 2136 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 4062 13812 4068 13864
rect 4120 13812 4126 13864
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 5626 13852 5632 13864
rect 5583 13824 5632 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9324 13852 9352 14019
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 10284 14028 11437 14056
rect 10284 14016 10290 14028
rect 11425 14025 11437 14028
rect 11471 14056 11483 14059
rect 11790 14056 11796 14068
rect 11471 14028 11796 14056
rect 11471 14025 11483 14028
rect 11425 14019 11483 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 18414 14056 18420 14068
rect 17727 14028 18420 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14056 20867 14059
rect 22186 14056 22192 14068
rect 20855 14028 22192 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 10686 13988 10692 14000
rect 10647 13960 10692 13988
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 11330 13988 11336 14000
rect 11195 13960 11336 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 11330 13948 11336 13960
rect 11388 13988 11394 14000
rect 13725 13991 13783 13997
rect 13725 13988 13737 13991
rect 11388 13960 13737 13988
rect 11388 13948 11394 13960
rect 13725 13957 13737 13960
rect 13771 13957 13783 13991
rect 13725 13951 13783 13957
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 15896 13960 16804 13988
rect 15896 13948 15902 13960
rect 9674 13920 9680 13932
rect 9635 13892 9680 13920
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 11882 13920 11888 13932
rect 9784 13892 11888 13920
rect 9784 13861 9812 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15930 13920 15936 13932
rect 14875 13892 15936 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16666 13920 16672 13932
rect 16500 13892 16672 13920
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9272 13824 9781 13852
rect 9272 13812 9278 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12768 13824 12817 13852
rect 12768 13812 12774 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12894 13812 12900 13864
rect 12952 13852 12958 13864
rect 13354 13852 13360 13864
rect 12952 13824 12997 13852
rect 13315 13824 13360 13852
rect 12952 13812 12958 13824
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 13538 13852 13544 13864
rect 13451 13824 13544 13852
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13852 16175 13855
rect 16163 13824 16197 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13784 2467 13787
rect 2958 13784 2964 13796
rect 2455 13756 2964 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 4706 13784 4712 13796
rect 4667 13756 4712 13784
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 6457 13787 6515 13793
rect 6457 13753 6469 13787
rect 6503 13784 6515 13787
rect 7282 13784 7288 13796
rect 6503 13756 7288 13784
rect 6503 13753 6515 13756
rect 6457 13747 6515 13753
rect 7282 13744 7288 13756
rect 7340 13744 7346 13796
rect 7926 13744 7932 13796
rect 7984 13744 7990 13796
rect 12069 13787 12127 13793
rect 12069 13753 12081 13787
rect 12115 13784 12127 13787
rect 13556 13784 13584 13812
rect 12115 13756 13584 13784
rect 16132 13784 16160 13815
rect 16390 13812 16396 13864
rect 16448 13852 16454 13864
rect 16500 13861 16528 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 16448 13824 16497 13852
rect 16448 13812 16454 13824
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 16577 13855 16635 13861
rect 16577 13821 16589 13855
rect 16623 13852 16635 13855
rect 16776 13852 16804 13960
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 20898 13988 20904 14000
rect 19484 13960 20904 13988
rect 19484 13948 19490 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 22465 13991 22523 13997
rect 22465 13988 22477 13991
rect 21416 13960 22477 13988
rect 21416 13948 21422 13960
rect 22465 13957 22477 13960
rect 22511 13988 22523 13991
rect 22922 13988 22928 14000
rect 22511 13960 22928 13988
rect 22511 13957 22523 13960
rect 22465 13951 22523 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 18831 13892 19533 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19521 13889 19533 13892
rect 19567 13920 19579 13923
rect 19978 13920 19984 13932
rect 19567 13892 19984 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20088 13892 21097 13920
rect 20088 13864 20116 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 21085 13883 21143 13889
rect 21652 13892 22845 13920
rect 16623 13824 16804 13852
rect 18417 13855 18475 13861
rect 16623 13821 16635 13824
rect 16577 13815 16635 13821
rect 18417 13821 18429 13855
rect 18463 13852 18475 13855
rect 19150 13852 19156 13864
rect 18463 13824 19156 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 20070 13852 20076 13864
rect 19983 13824 20076 13852
rect 19705 13815 19763 13821
rect 16942 13784 16948 13796
rect 16132 13756 16948 13784
rect 12115 13753 12127 13756
rect 12069 13747 12127 13753
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 17313 13787 17371 13793
rect 17313 13753 17325 13787
rect 17359 13784 17371 13787
rect 18782 13784 18788 13796
rect 17359 13756 18788 13784
rect 17359 13753 17371 13756
rect 17313 13747 17371 13753
rect 18782 13744 18788 13756
rect 18840 13784 18846 13796
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18840 13756 19073 13784
rect 18840 13744 18846 13756
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 19242 13744 19248 13796
rect 19300 13784 19306 13796
rect 19720 13784 19748 13815
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 20254 13852 20260 13864
rect 20215 13824 20260 13852
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 21652 13861 21680 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21637 13815 21695 13821
rect 21652 13784 21680 13815
rect 19300 13756 21680 13784
rect 19300 13744 19306 13756
rect 15194 13716 15200 13728
rect 15155 13688 15200 13716
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 15562 13716 15568 13728
rect 15523 13688 15568 13716
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20070 13716 20076 13728
rect 19392 13688 20076 13716
rect 19392 13676 19398 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 22094 13716 22100 13728
rect 22055 13688 22100 13716
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 1104 13626 24656 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 24656 13626
rect 1104 13552 24656 13574
rect 2590 13512 2596 13524
rect 2551 13484 2596 13512
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 3016 13484 5396 13512
rect 3016 13472 3022 13484
rect 3237 13447 3295 13453
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 4062 13444 4068 13456
rect 3283 13416 4068 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 4632 13416 5304 13444
rect 5368 13416 5396 13484
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 7340 13484 8309 13512
rect 7340 13472 7346 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 8297 13475 8355 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 13354 13512 13360 13524
rect 12575 13484 13360 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 14182 13512 14188 13524
rect 14143 13484 14188 13512
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15746 13512 15752 13524
rect 15252 13484 15752 13512
rect 15252 13472 15258 13484
rect 15746 13472 15752 13484
rect 15804 13512 15810 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 15804 13484 16681 13512
rect 15804 13472 15810 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 17129 13515 17187 13521
rect 17129 13512 17141 13515
rect 17000 13484 17141 13512
rect 17000 13472 17006 13484
rect 17129 13481 17141 13484
rect 17175 13481 17187 13515
rect 19150 13512 19156 13524
rect 19111 13484 19156 13512
rect 17129 13475 17187 13481
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13512 19487 13515
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19475 13484 19809 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 6825 13447 6883 13453
rect 4632 13388 4660 13416
rect 2774 13376 2780 13388
rect 2735 13348 2780 13376
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4614 13376 4620 13388
rect 4575 13348 4620 13376
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5276 13376 5304 13416
rect 6825 13413 6837 13447
rect 6871 13444 6883 13447
rect 7650 13444 7656 13456
rect 6871 13416 7656 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 7650 13404 7656 13416
rect 7708 13444 7714 13456
rect 7926 13444 7932 13456
rect 7708 13416 7932 13444
rect 7708 13404 7714 13416
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 10137 13447 10195 13453
rect 10137 13444 10149 13447
rect 9824 13416 10149 13444
rect 9824 13404 9830 13416
rect 10137 13413 10149 13416
rect 10183 13413 10195 13447
rect 10137 13407 10195 13413
rect 10594 13404 10600 13456
rect 10652 13404 10658 13456
rect 11882 13444 11888 13456
rect 11843 13416 11888 13444
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 13173 13447 13231 13453
rect 13173 13444 13185 13447
rect 12768 13416 13185 13444
rect 12768 13404 12774 13416
rect 13173 13413 13185 13416
rect 13219 13413 13231 13447
rect 13173 13407 13231 13413
rect 14921 13447 14979 13453
rect 14921 13413 14933 13447
rect 14967 13444 14979 13447
rect 17773 13447 17831 13453
rect 14967 13416 16252 13444
rect 14967 13413 14979 13416
rect 14921 13407 14979 13413
rect 7098 13376 7104 13388
rect 5276 13348 7104 13376
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7248 13348 7297 13376
rect 7248 13336 7254 13348
rect 7285 13345 7297 13348
rect 7331 13376 7343 13379
rect 7466 13376 7472 13388
rect 7331 13348 7472 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 7837 13379 7895 13385
rect 7837 13376 7849 13379
rect 7800 13348 7849 13376
rect 7800 13336 7806 13348
rect 7837 13345 7849 13348
rect 7883 13345 7895 13379
rect 8018 13376 8024 13388
rect 7979 13348 8024 13376
rect 7837 13339 7895 13345
rect 8018 13336 8024 13348
rect 8076 13336 8082 13388
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15620 13348 15669 13376
rect 15620 13336 15626 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16224 13385 16252 13416
rect 17773 13413 17785 13447
rect 17819 13444 17831 13447
rect 19242 13444 19248 13456
rect 17819 13416 19248 13444
rect 17819 13413 17831 13416
rect 17773 13407 17831 13413
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 20533 13447 20591 13453
rect 20533 13413 20545 13447
rect 20579 13444 20591 13447
rect 21358 13444 21364 13456
rect 20579 13416 21364 13444
rect 20579 13413 20591 13416
rect 20533 13407 20591 13413
rect 21358 13404 21364 13416
rect 21416 13444 21422 13456
rect 21416 13416 21772 13444
rect 21416 13404 21422 13416
rect 16117 13379 16175 13385
rect 16117 13376 16129 13379
rect 15896 13348 16129 13376
rect 15896 13336 15902 13348
rect 16117 13345 16129 13348
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16209 13379 16267 13385
rect 16209 13345 16221 13379
rect 16255 13376 16267 13379
rect 16758 13376 16764 13388
rect 16255 13348 16764 13376
rect 16255 13345 16267 13348
rect 16209 13339 16267 13345
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 18414 13376 18420 13388
rect 17920 13348 18420 13376
rect 17920 13336 17926 13348
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 21542 13376 21548 13388
rect 21503 13348 21548 13376
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 21744 13385 21772 13416
rect 22094 13404 22100 13456
rect 22152 13404 22158 13456
rect 21729 13379 21787 13385
rect 21729 13345 21741 13379
rect 21775 13345 21787 13379
rect 21729 13339 21787 13345
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 7208 13240 7236 13336
rect 9858 13308 9864 13320
rect 9819 13280 9864 13308
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 5224 13212 7236 13240
rect 15488 13240 15516 13271
rect 15654 13240 15660 13252
rect 15488 13212 15660 13240
rect 5224 13200 5230 13212
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 2188 13144 3525 13172
rect 2188 13132 2194 13144
rect 3513 13141 3525 13144
rect 3559 13141 3571 13175
rect 3513 13135 3571 13141
rect 3602 13132 3608 13184
rect 3660 13172 3666 13184
rect 7558 13172 7564 13184
rect 3660 13144 7564 13172
rect 3660 13132 3666 13144
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18601 13175 18659 13181
rect 18601 13172 18613 13175
rect 18187 13144 18613 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18601 13141 18613 13144
rect 18647 13172 18659 13175
rect 18966 13172 18972 13184
rect 18647 13144 18972 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 1104 13082 24656 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 24656 13082
rect 1104 13008 24656 13030
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 2740 12940 3157 12968
rect 2740 12928 2746 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3145 12931 3203 12937
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4614 12968 4620 12980
rect 4479 12940 4620 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 1596 12696 1624 12727
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 3160 12764 3188 12931
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 5166 12968 5172 12980
rect 4847 12940 5172 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5534 12968 5540 12980
rect 5495 12940 5540 12968
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 8202 12968 8208 12980
rect 7156 12940 8208 12968
rect 7156 12928 7162 12940
rect 8202 12928 8208 12940
rect 8260 12968 8266 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 8260 12940 8309 12968
rect 8260 12928 8266 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 8297 12931 8355 12937
rect 10137 12971 10195 12977
rect 10137 12937 10149 12971
rect 10183 12968 10195 12971
rect 10594 12968 10600 12980
rect 10183 12940 10600 12968
rect 10183 12937 10195 12940
rect 10137 12931 10195 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 15896 12940 16405 12968
rect 15896 12928 15902 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 16758 12968 16764 12980
rect 16719 12940 16764 12968
rect 16393 12931 16451 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17218 12968 17224 12980
rect 17179 12940 17224 12968
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 3421 12903 3479 12909
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 4706 12900 4712 12912
rect 3467 12872 4712 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 7466 12860 7472 12912
rect 7524 12900 7530 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 7524 12872 8677 12900
rect 7524 12860 7530 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 8665 12863 8723 12869
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6503 12804 7297 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 7285 12801 7297 12804
rect 7331 12832 7343 12835
rect 8018 12832 8024 12844
rect 7331 12804 8024 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 20257 12835 20315 12841
rect 20257 12832 20269 12835
rect 19300 12804 20269 12832
rect 19300 12792 19306 12804
rect 20257 12801 20269 12804
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 5350 12764 5356 12776
rect 1728 12736 1773 12764
rect 3160 12736 4154 12764
rect 5311 12736 5356 12764
rect 1728 12724 1734 12736
rect 2869 12699 2927 12705
rect 2869 12696 2881 12699
rect 1596 12668 2881 12696
rect 2869 12665 2881 12668
rect 2915 12696 2927 12699
rect 3602 12696 3608 12708
rect 2915 12668 3608 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 4126 12696 4154 12736
rect 5350 12724 5356 12736
rect 5408 12764 5414 12776
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 5408 12736 5825 12764
rect 5408 12724 5414 12736
rect 5813 12733 5825 12736
rect 5859 12733 5871 12767
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 5813 12727 5871 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 14366 12764 14372 12776
rect 13955 12736 14372 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 14516 12736 15117 12764
rect 14516 12724 14522 12736
rect 15105 12733 15117 12736
rect 15151 12764 15163 12767
rect 15562 12764 15568 12776
rect 15151 12736 15568 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 15562 12724 15568 12736
rect 15620 12764 15626 12776
rect 16298 12764 16304 12776
rect 15620 12736 16304 12764
rect 15620 12724 15626 12736
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 18230 12764 18236 12776
rect 17276 12736 18236 12764
rect 17276 12724 17282 12736
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12764 20775 12767
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20763 12736 21005 12764
rect 20763 12733 20775 12736
rect 20717 12727 20775 12733
rect 20993 12733 21005 12736
rect 21039 12764 21051 12767
rect 21450 12764 21456 12776
rect 21039 12736 21456 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 21729 12767 21787 12773
rect 21729 12733 21741 12767
rect 21775 12764 21787 12767
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21775 12736 22109 12764
rect 21775 12733 21787 12736
rect 21729 12727 21787 12733
rect 22097 12733 22109 12736
rect 22143 12764 22155 12767
rect 22462 12764 22468 12776
rect 22143 12736 22468 12764
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 22462 12724 22468 12736
rect 22520 12764 22526 12776
rect 23382 12764 23388 12776
rect 22520 12736 23388 12764
rect 22520 12724 22526 12736
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 6914 12696 6920 12708
rect 4126 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12696 6978 12708
rect 9309 12699 9367 12705
rect 9309 12696 9321 12699
rect 6972 12668 9321 12696
rect 6972 12656 6978 12668
rect 9309 12665 9321 12668
rect 9355 12696 9367 12699
rect 9858 12696 9864 12708
rect 9355 12668 9864 12696
rect 9355 12665 9367 12668
rect 9309 12659 9367 12665
rect 9858 12656 9864 12668
rect 9916 12696 9922 12708
rect 11149 12699 11207 12705
rect 9916 12668 10732 12696
rect 9916 12656 9922 12668
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3421 12631 3479 12637
rect 3421 12628 3433 12631
rect 2832 12600 3433 12628
rect 2832 12588 2838 12600
rect 3421 12597 3433 12600
rect 3467 12628 3479 12631
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 3467 12600 3525 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 9766 12628 9772 12640
rect 9727 12600 9772 12628
rect 3513 12591 3571 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10594 12628 10600 12640
rect 10551 12600 10600 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10704 12628 10732 12668
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 11977 12699 12035 12705
rect 11977 12696 11989 12699
rect 11195 12668 11989 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 11977 12665 11989 12668
rect 12023 12696 12035 12699
rect 12618 12696 12624 12708
rect 12023 12668 12624 12696
rect 12023 12665 12035 12668
rect 11977 12659 12035 12665
rect 12618 12656 12624 12668
rect 12676 12696 12682 12708
rect 12713 12699 12771 12705
rect 12713 12696 12725 12699
rect 12676 12668 12725 12696
rect 12676 12656 12682 12668
rect 12713 12665 12725 12668
rect 12759 12665 12771 12699
rect 12713 12659 12771 12665
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 14918 12696 14924 12708
rect 13127 12668 14924 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 15470 12656 15476 12708
rect 15528 12656 15534 12708
rect 17681 12699 17739 12705
rect 17681 12665 17693 12699
rect 17727 12696 17739 12699
rect 18506 12696 18512 12708
rect 17727 12668 18512 12696
rect 17727 12665 17739 12668
rect 17681 12659 17739 12665
rect 18506 12656 18512 12668
rect 18564 12656 18570 12708
rect 18966 12656 18972 12708
rect 19024 12656 19030 12708
rect 22002 12696 22008 12708
rect 21963 12668 22008 12696
rect 22002 12656 22008 12668
rect 22060 12656 22066 12708
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 10704 12600 11253 12628
rect 11241 12597 11253 12600
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21542 12628 21548 12640
rect 21223 12600 21548 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21542 12588 21548 12600
rect 21600 12628 21606 12640
rect 21726 12628 21732 12640
rect 21600 12600 21732 12628
rect 21600 12588 21606 12600
rect 21726 12588 21732 12600
rect 21784 12588 21790 12640
rect 1104 12538 24656 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 24656 12538
rect 1104 12464 24656 12486
rect 2501 12427 2559 12433
rect 2501 12393 2513 12427
rect 2547 12424 2559 12427
rect 2590 12424 2596 12436
rect 2547 12396 2596 12424
rect 2547 12393 2559 12396
rect 2501 12387 2559 12393
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 2774 12424 2780 12436
rect 2735 12396 2780 12424
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 5350 12424 5356 12436
rect 5311 12396 5356 12424
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7742 12424 7748 12436
rect 7703 12396 7748 12424
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8202 12424 8208 12436
rect 8163 12396 8208 12424
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 12618 12424 12624 12436
rect 9824 12396 11468 12424
rect 12579 12396 12624 12424
rect 9824 12384 9830 12396
rect 1118 12248 1124 12300
rect 1176 12288 1182 12300
rect 1670 12288 1676 12300
rect 1176 12260 1676 12288
rect 1176 12248 1182 12260
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5074 12288 5080 12300
rect 4939 12260 5080 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5074 12248 5080 12260
rect 5132 12288 5138 12300
rect 5368 12288 5396 12384
rect 11440 12328 11468 12396
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 14458 12424 14464 12436
rect 14419 12396 14464 12424
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 15470 12424 15476 12436
rect 15431 12396 15476 12424
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16298 12424 16304 12436
rect 16259 12396 16304 12424
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 17276 12396 17693 12424
rect 17276 12384 17282 12396
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 19981 12427 20039 12433
rect 19981 12424 19993 12427
rect 18932 12396 19993 12424
rect 18932 12384 18938 12396
rect 19981 12393 19993 12396
rect 20027 12393 20039 12427
rect 19981 12387 20039 12393
rect 20533 12359 20591 12365
rect 20533 12325 20545 12359
rect 20579 12356 20591 12359
rect 21726 12356 21732 12368
rect 20579 12328 21732 12356
rect 20579 12325 20591 12328
rect 20533 12319 20591 12325
rect 21726 12316 21732 12328
rect 21784 12316 21790 12368
rect 22094 12316 22100 12368
rect 22152 12316 22158 12368
rect 23382 12356 23388 12368
rect 23343 12328 23388 12356
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 8018 12288 8024 12300
rect 5132 12260 5396 12288
rect 7979 12260 8024 12288
rect 5132 12248 5138 12260
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10183 12260 10517 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1544 12192 1593 12220
rect 1544 12180 1550 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 1581 12183 1639 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 4798 12152 4804 12164
rect 3160 12124 4804 12152
rect 3160 12096 3188 12124
rect 4798 12112 4804 12124
rect 4856 12152 4862 12164
rect 5626 12152 5632 12164
rect 4856 12124 5632 12152
rect 4856 12112 4862 12124
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 10520 12152 10548 12251
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 10652 12260 11345 12288
rect 10652 12248 10658 12260
rect 11333 12257 11345 12260
rect 11379 12288 11391 12291
rect 12710 12288 12716 12300
rect 11379 12260 12716 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 13906 12288 13912 12300
rect 13219 12260 13912 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 13906 12248 13912 12260
rect 13964 12288 13970 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13964 12260 14013 12288
rect 13964 12248 13970 12260
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 15930 12288 15936 12300
rect 15887 12260 15936 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 15930 12248 15936 12260
rect 15988 12288 15994 12300
rect 18414 12288 18420 12300
rect 15988 12260 18420 12288
rect 15988 12248 15994 12260
rect 18414 12248 18420 12260
rect 18472 12288 18478 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18472 12260 18797 12288
rect 18472 12248 18478 12260
rect 18785 12257 18797 12260
rect 18831 12288 18843 12291
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 18831 12260 19257 12288
rect 18831 12257 18843 12260
rect 18785 12251 18843 12257
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 20622 12288 20628 12300
rect 19843 12260 20628 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21361 12291 21419 12297
rect 21361 12288 21373 12291
rect 21140 12260 21373 12288
rect 21140 12248 21146 12260
rect 21361 12257 21373 12260
rect 21407 12257 21419 12291
rect 21361 12251 21419 12257
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 13630 12220 13636 12232
rect 12584 12192 13636 12220
rect 12584 12180 12590 12192
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 21634 12220 21640 12232
rect 21595 12192 21640 12220
rect 21634 12180 21640 12192
rect 21692 12180 21698 12232
rect 12802 12152 12808 12164
rect 10520 12124 12808 12152
rect 12802 12112 12808 12124
rect 12860 12152 12866 12164
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 12860 12124 13369 12152
rect 12860 12112 12866 12124
rect 13357 12121 13369 12124
rect 13403 12121 13415 12155
rect 13357 12115 13415 12121
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18187 12124 19012 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18984 12096 19012 12124
rect 3142 12084 3148 12096
rect 3103 12056 3148 12084
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3602 12084 3608 12096
rect 3563 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 5040 12056 5089 12084
rect 5040 12044 5046 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14424 12056 14933 12084
rect 14424 12044 14430 12056
rect 14921 12053 14933 12056
rect 14967 12084 14979 12087
rect 15654 12084 15660 12096
rect 14967 12056 15660 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16022 12084 16028 12096
rect 15983 12056 16028 12084
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 18966 12084 18972 12096
rect 18927 12056 18972 12084
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 1104 11994 24656 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 24656 11994
rect 1104 11920 24656 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 10505 11883 10563 11889
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 10870 11880 10876 11892
rect 10551 11852 10876 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 1486 11772 1492 11824
rect 1544 11812 1550 11824
rect 9217 11815 9275 11821
rect 9217 11812 9229 11815
rect 1544 11784 3740 11812
rect 1544 11772 1550 11784
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 3712 11744 3740 11784
rect 5460 11784 9229 11812
rect 5460 11744 5488 11784
rect 9217 11781 9229 11784
rect 9263 11812 9275 11815
rect 9493 11815 9551 11821
rect 9493 11812 9505 11815
rect 9263 11784 9505 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 9493 11781 9505 11784
rect 9539 11781 9551 11815
rect 9493 11775 9551 11781
rect 5626 11744 5632 11756
rect 3712 11716 5488 11744
rect 5587 11716 5632 11744
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8018 11744 8024 11756
rect 7975 11716 8024 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8018 11704 8024 11716
rect 8076 11744 8082 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 8076 11716 10241 11744
rect 8076 11704 8082 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3142 11676 3148 11688
rect 2731 11648 3148 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 4982 11636 4988 11688
rect 5040 11636 5046 11688
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9582 11676 9588 11688
rect 9539 11648 9588 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 3329 11611 3387 11617
rect 3329 11577 3341 11611
rect 3375 11608 3387 11611
rect 3878 11608 3884 11620
rect 3375 11580 3884 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 8588 11608 8616 11639
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10520 11676 10548 11843
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 12805 11883 12863 11889
rect 12805 11880 12817 11883
rect 12584 11852 12817 11880
rect 12584 11840 12590 11852
rect 12805 11849 12817 11852
rect 12851 11849 12863 11883
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 12805 11843 12863 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14090 11812 14096 11824
rect 13096 11784 14096 11812
rect 10962 11676 10968 11688
rect 9723 11648 10548 11676
rect 10923 11648 10968 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11103 11648 11928 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 8343 11580 10149 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 10229 11611 10287 11617
rect 10229 11577 10241 11611
rect 10275 11608 10287 11611
rect 11517 11611 11575 11617
rect 11517 11608 11529 11611
rect 10275 11580 11529 11608
rect 10275 11577 10287 11580
rect 10229 11571 10287 11577
rect 11517 11577 11529 11580
rect 11563 11577 11575 11611
rect 11517 11571 11575 11577
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 11900 11549 11928 11648
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 13096 11685 13124 11784
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 21085 11815 21143 11821
rect 21085 11781 21097 11815
rect 21131 11812 21143 11815
rect 21634 11812 21640 11824
rect 21131 11784 21640 11812
rect 21131 11781 21143 11784
rect 21085 11775 21143 11781
rect 21634 11772 21640 11784
rect 21692 11812 21698 11824
rect 22465 11815 22523 11821
rect 22465 11812 22477 11815
rect 21692 11784 22477 11812
rect 21692 11772 21698 11784
rect 22465 11781 22477 11784
rect 22511 11781 22523 11815
rect 22465 11775 22523 11781
rect 13630 11744 13636 11756
rect 13591 11716 13636 11744
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 14918 11704 14924 11756
rect 14976 11744 14982 11756
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14976 11716 15025 11744
rect 14976 11704 14982 11716
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15378 11744 15384 11756
rect 15335 11716 15384 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 18230 11744 18236 11756
rect 18191 11716 18236 11744
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12492 11648 12633 11676
rect 12492 11636 12498 11648
rect 12621 11645 12633 11648
rect 12667 11676 12679 11679
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 12667 11648 13093 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 13081 11645 13093 11648
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 7156 11512 8769 11540
rect 7156 11500 7162 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12066 11540 12072 11552
rect 11931 11512 12072 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 13740 11540 13768 11639
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 21545 11679 21603 11685
rect 21545 11676 21557 11679
rect 21416 11648 21557 11676
rect 21416 11636 21422 11648
rect 21545 11645 21557 11648
rect 21591 11645 21603 11679
rect 21545 11639 21603 11645
rect 21637 11679 21695 11685
rect 21637 11645 21649 11679
rect 21683 11676 21695 11679
rect 21726 11676 21732 11688
rect 21683 11648 21732 11676
rect 21683 11645 21695 11648
rect 21637 11639 21695 11645
rect 21726 11636 21732 11648
rect 21784 11636 21790 11688
rect 22002 11676 22008 11688
rect 21963 11648 22008 11676
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11676 22155 11679
rect 22186 11676 22192 11688
rect 22143 11648 22192 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 16022 11568 16028 11620
rect 16080 11568 16086 11620
rect 16850 11568 16856 11620
rect 16908 11608 16914 11620
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 16908 11580 17049 11608
rect 16908 11568 16914 11580
rect 17037 11577 17049 11580
rect 17083 11577 17095 11611
rect 17037 11571 17095 11577
rect 17681 11611 17739 11617
rect 17681 11577 17693 11611
rect 17727 11608 17739 11611
rect 18509 11611 18567 11617
rect 18509 11608 18521 11611
rect 17727 11580 18521 11608
rect 17727 11577 17739 11580
rect 17681 11571 17739 11577
rect 18509 11577 18521 11580
rect 18555 11608 18567 11611
rect 18598 11608 18604 11620
rect 18555 11580 18604 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 18598 11568 18604 11580
rect 18656 11568 18662 11620
rect 18966 11568 18972 11620
rect 19024 11568 19030 11620
rect 20257 11611 20315 11617
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 20346 11608 20352 11620
rect 20303 11580 20352 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 13740 11512 14565 11540
rect 14553 11509 14565 11512
rect 14599 11540 14611 11543
rect 15102 11540 15108 11552
rect 14599 11512 15108 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 20622 11540 20628 11552
rect 20583 11512 20628 11540
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 21744 11540 21772 11636
rect 22020 11608 22048 11636
rect 23017 11611 23075 11617
rect 23017 11608 23029 11611
rect 22020 11580 23029 11608
rect 23017 11577 23029 11580
rect 23063 11577 23075 11611
rect 23017 11571 23075 11577
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 21744 11512 23857 11540
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 1104 11450 24656 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 24656 11450
rect 1104 11376 24656 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2188 11308 2421 11336
rect 2188 11296 2194 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 3936 11308 5764 11336
rect 3936 11296 3942 11308
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 2148 11200 2176 11296
rect 3697 11271 3755 11277
rect 3697 11237 3709 11271
rect 3743 11268 3755 11271
rect 4982 11268 4988 11280
rect 3743 11240 4988 11268
rect 3743 11237 3755 11240
rect 3697 11231 3755 11237
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 5736 11240 5764 11308
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 10045 11339 10103 11345
rect 10045 11336 10057 11339
rect 7616 11308 10057 11336
rect 7616 11296 7622 11308
rect 10045 11305 10057 11308
rect 10091 11336 10103 11339
rect 10413 11339 10471 11345
rect 10413 11336 10425 11339
rect 10091 11308 10425 11336
rect 10091 11305 10103 11308
rect 10045 11299 10103 11305
rect 10413 11305 10425 11308
rect 10459 11336 10471 11339
rect 10962 11336 10968 11348
rect 10459 11308 10968 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 14921 11339 14979 11345
rect 14921 11305 14933 11339
rect 14967 11336 14979 11339
rect 16022 11336 16028 11348
rect 14967 11308 16028 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 20956 11308 21281 11336
rect 20956 11296 20962 11308
rect 21269 11305 21281 11308
rect 21315 11305 21327 11339
rect 21269 11299 21327 11305
rect 21637 11339 21695 11345
rect 21637 11305 21649 11339
rect 21683 11336 21695 11339
rect 22094 11336 22100 11348
rect 21683 11308 22100 11336
rect 21683 11305 21695 11308
rect 21637 11299 21695 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 12434 11268 12440 11280
rect 9876 11240 12440 11268
rect 9876 11212 9904 11240
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 12529 11271 12587 11277
rect 12529 11237 12541 11271
rect 12575 11268 12587 11271
rect 12618 11268 12624 11280
rect 12575 11240 12624 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 12618 11228 12624 11240
rect 12676 11268 12682 11280
rect 13449 11271 13507 11277
rect 13449 11268 13461 11271
rect 12676 11240 13461 11268
rect 12676 11228 12682 11240
rect 13449 11237 13461 11240
rect 13495 11237 13507 11271
rect 15930 11268 15936 11280
rect 15891 11240 15936 11268
rect 13449 11231 13507 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 16853 11271 16911 11277
rect 16853 11237 16865 11271
rect 16899 11268 16911 11271
rect 16899 11240 18092 11268
rect 16899 11237 16911 11240
rect 16853 11231 16911 11237
rect 5626 11200 5632 11212
rect 1627 11172 2176 11200
rect 5587 11172 5632 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6362 11200 6368 11212
rect 6135 11172 6368 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6362 11160 6368 11172
rect 6420 11200 6426 11212
rect 7098 11200 7104 11212
rect 6420 11172 7104 11200
rect 6420 11160 6426 11172
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 7524 11172 7573 11200
rect 7524 11160 7530 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 9858 11200 9864 11212
rect 9819 11172 9864 11200
rect 7561 11163 7619 11169
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 14918 11200 14924 11212
rect 14599 11172 14924 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7742 11132 7748 11144
rect 7055 11104 7748 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 10796 11132 10824 11163
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15746 11200 15752 11212
rect 15519 11172 15752 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 18064 11209 18092 11240
rect 18506 11228 18512 11280
rect 18564 11228 18570 11280
rect 20533 11271 20591 11277
rect 20533 11237 20545 11271
rect 20579 11268 20591 11271
rect 22186 11268 22192 11280
rect 20579 11240 22192 11268
rect 20579 11237 20591 11240
rect 20533 11231 20591 11237
rect 22186 11228 22192 11240
rect 22244 11268 22250 11280
rect 22244 11240 23060 11268
rect 22244 11228 22250 11240
rect 23032 11212 23060 11240
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18414 11200 18420 11212
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 10870 11132 10876 11144
rect 10796 11104 10876 11132
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 1765 11067 1823 11073
rect 1765 11033 1777 11067
rect 1811 11064 1823 11067
rect 1854 11064 1860 11076
rect 1811 11036 1860 11064
rect 1811 11033 1823 11036
rect 1765 11027 1823 11033
rect 1854 11024 1860 11036
rect 1912 11064 1918 11076
rect 13630 11064 13636 11076
rect 1912 11036 2176 11064
rect 13591 11036 13636 11064
rect 1912 11024 1918 11036
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 2041 10999 2099 11005
rect 2041 10996 2053 10999
rect 1544 10968 2053 10996
rect 1544 10956 1550 10968
rect 2041 10965 2053 10968
rect 2087 10965 2099 10999
rect 2148 10996 2176 11036
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 15654 11064 15660 11076
rect 15615 11036 15660 11064
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 17420 11064 17448 11163
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 21085 11203 21143 11209
rect 21085 11169 21097 11203
rect 21131 11200 21143 11203
rect 21266 11200 21272 11212
rect 21131 11172 21272 11200
rect 21131 11169 21143 11172
rect 21085 11163 21143 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 22005 11203 22063 11209
rect 22005 11200 22017 11203
rect 21416 11172 22017 11200
rect 21416 11160 21422 11172
rect 22005 11169 22017 11172
rect 22051 11169 22063 11203
rect 22462 11200 22468 11212
rect 22423 11172 22468 11200
rect 22005 11163 22063 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22646 11200 22652 11212
rect 22607 11172 22652 11200
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 23014 11200 23020 11212
rect 22927 11172 23020 11200
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 18506 11064 18512 11076
rect 17420 11036 18512 11064
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 20165 11067 20223 11073
rect 20165 11033 20177 11067
rect 20211 11064 20223 11067
rect 21082 11064 21088 11076
rect 20211 11036 21088 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 22002 11024 22008 11076
rect 22060 11064 22066 11076
rect 22940 11064 22968 11095
rect 22060 11036 22968 11064
rect 22060 11024 22066 11036
rect 2866 10996 2872 11008
rect 2148 10968 2872 10996
rect 2041 10959 2099 10965
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 3237 10999 3295 11005
rect 3237 10965 3249 10999
rect 3283 10996 3295 10999
rect 3602 10996 3608 11008
rect 3283 10968 3608 10996
rect 3283 10965 3295 10968
rect 3237 10959 3295 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4249 10999 4307 11005
rect 4249 10996 4261 10999
rect 4028 10968 4261 10996
rect 4028 10956 4034 10968
rect 4249 10965 4261 10968
rect 4295 10965 4307 10999
rect 4249 10959 4307 10965
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7064 10968 7757 10996
rect 7064 10956 7070 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 1104 10906 24656 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 24656 10906
rect 1104 10832 24656 10854
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5684 10764 6009 10792
rect 5684 10752 5690 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 10870 10792 10876 10804
rect 10827 10764 10876 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12618 10792 12624 10804
rect 11931 10764 12624 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4028 10628 5089 10656
rect 4028 10616 4034 10628
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6972 10628 7021 10656
rect 6972 10616 6978 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9858 10656 9864 10668
rect 9447 10628 9864 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9858 10616 9864 10628
rect 9916 10656 9922 10668
rect 10226 10656 10232 10668
rect 9916 10628 10232 10656
rect 9916 10616 9922 10628
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 1854 10588 1860 10600
rect 1815 10560 1860 10588
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2038 10548 2044 10600
rect 2096 10588 2102 10600
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 2096 10560 2513 10588
rect 2096 10548 2102 10560
rect 2501 10557 2513 10560
rect 2547 10588 2559 10591
rect 3881 10591 3939 10597
rect 2547 10560 3648 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3620 10532 3648 10560
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 4062 10588 4068 10600
rect 3927 10560 4068 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 4062 10548 4068 10560
rect 4120 10588 4126 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4120 10560 4629 10588
rect 4120 10548 4126 10560
rect 4617 10557 4629 10560
rect 4663 10588 4675 10591
rect 4706 10588 4712 10600
rect 4663 10560 4712 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 5169 10591 5227 10597
rect 4856 10560 4901 10588
rect 4856 10548 4862 10560
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 9674 10588 9680 10600
rect 9587 10560 9680 10588
rect 5169 10551 5227 10557
rect 3510 10520 3516 10532
rect 3471 10492 3516 10520
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 4157 10523 4215 10529
rect 4157 10520 4169 10523
rect 3660 10492 4169 10520
rect 3660 10480 3666 10492
rect 4157 10489 4169 10492
rect 4203 10489 4215 10523
rect 4157 10483 4215 10489
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 4614 10452 4620 10464
rect 2556 10424 4620 10452
rect 2556 10412 2562 10424
rect 4614 10412 4620 10424
rect 4672 10452 4678 10464
rect 5184 10452 5212 10551
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 11149 10591 11207 10597
rect 9732 10560 10272 10588
rect 9732 10548 9738 10560
rect 6457 10523 6515 10529
rect 6457 10489 6469 10523
rect 6503 10520 6515 10523
rect 7282 10520 7288 10532
rect 6503 10492 7288 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 7742 10480 7748 10532
rect 7800 10480 7806 10532
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10489 9091 10523
rect 9033 10483 9091 10489
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 4672 10424 5641 10452
rect 4672 10412 4678 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 9048 10452 9076 10483
rect 9858 10452 9864 10464
rect 7524 10424 9076 10452
rect 9819 10424 9864 10452
rect 7524 10412 7530 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10244 10461 10272 10560
rect 11149 10557 11161 10591
rect 11195 10588 11207 10591
rect 11900 10588 11928 10755
rect 12618 10752 12624 10764
rect 12676 10792 12682 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 12676 10764 13461 10792
rect 12676 10752 12682 10764
rect 13449 10761 13461 10764
rect 13495 10761 13507 10795
rect 14090 10792 14096 10804
rect 14051 10764 14096 10792
rect 13449 10755 13507 10761
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14734 10792 14740 10804
rect 14695 10764 14740 10792
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 22005 10795 22063 10801
rect 22005 10761 22017 10795
rect 22051 10792 22063 10795
rect 22094 10792 22100 10804
rect 22051 10764 22100 10792
rect 22051 10761 22063 10764
rect 22005 10755 22063 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 22373 10795 22431 10801
rect 22373 10761 22385 10795
rect 22419 10792 22431 10795
rect 22462 10792 22468 10804
rect 22419 10764 22468 10792
rect 22419 10761 22431 10764
rect 22373 10755 22431 10761
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 14108 10656 14136 10752
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 19337 10727 19395 10733
rect 19337 10724 19349 10727
rect 18656 10696 19349 10724
rect 18656 10684 18662 10696
rect 19337 10693 19349 10696
rect 19383 10693 19395 10727
rect 19337 10687 19395 10693
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 14108 10628 14473 10656
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 22370 10656 22376 10668
rect 14461 10619 14519 10625
rect 21836 10628 22376 10656
rect 11195 10560 11928 10588
rect 12621 10591 12679 10597
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 13078 10588 13084 10600
rect 12667 10560 13084 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 15378 10588 15384 10600
rect 14599 10560 15384 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16850 10588 16856 10600
rect 16163 10560 16856 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 18969 10591 19027 10597
rect 18564 10560 18609 10588
rect 18564 10548 18570 10560
rect 18969 10557 18981 10591
rect 19015 10557 19027 10591
rect 19150 10588 19156 10600
rect 19063 10560 19156 10588
rect 18969 10551 19027 10557
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 17129 10523 17187 10529
rect 10376 10492 11284 10520
rect 10376 10480 10382 10492
rect 10229 10455 10287 10461
rect 10229 10421 10241 10455
rect 10275 10452 10287 10455
rect 10686 10452 10692 10464
rect 10275 10424 10692 10452
rect 10275 10421 10287 10424
rect 10229 10415 10287 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11256 10461 11284 10492
rect 17129 10489 17141 10523
rect 17175 10520 17187 10523
rect 18322 10520 18328 10532
rect 17175 10492 18328 10520
rect 17175 10489 17187 10492
rect 17129 10483 17187 10489
rect 18322 10480 18328 10492
rect 18380 10520 18386 10532
rect 18984 10520 19012 10551
rect 19150 10548 19156 10560
rect 19208 10588 19214 10600
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 19208 10560 20269 10588
rect 19208 10548 19214 10560
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 20346 10548 20352 10600
rect 20404 10588 20410 10600
rect 20404 10560 20497 10588
rect 20404 10548 20410 10560
rect 20530 10548 20536 10600
rect 20588 10588 20594 10600
rect 21836 10597 21864 10628
rect 22370 10616 22376 10628
rect 22428 10656 22434 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22428 10628 22661 10656
rect 22428 10616 22434 10628
rect 22649 10625 22661 10628
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 20588 10560 21833 10588
rect 20588 10548 20594 10560
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 21821 10551 21879 10557
rect 18380 10492 19012 10520
rect 18380 10480 18386 10492
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10421 11299 10455
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 11241 10415 11299 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 17681 10455 17739 10461
rect 17681 10421 17693 10455
rect 17727 10452 17739 10455
rect 17862 10452 17868 10464
rect 17727 10424 17868 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19889 10455 19947 10461
rect 19889 10452 19901 10455
rect 19484 10424 19901 10452
rect 19484 10412 19490 10424
rect 19889 10421 19901 10424
rect 19935 10452 19947 10455
rect 20364 10452 20392 10548
rect 22738 10480 22744 10532
rect 22796 10520 22802 10532
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 22796 10492 23857 10520
rect 22796 10480 22802 10492
rect 23845 10489 23857 10492
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 21266 10452 21272 10464
rect 19935 10424 20392 10452
rect 21227 10424 21272 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 21266 10412 21272 10424
rect 21324 10412 21330 10464
rect 1104 10362 24656 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 24656 10362
rect 1104 10288 24656 10310
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 3602 10248 3608 10260
rect 3559 10220 3608 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 4856 10220 5641 10248
rect 4856 10208 4862 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 5629 10211 5687 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 7800 10220 8493 10248
rect 7800 10208 7806 10220
rect 8481 10217 8493 10220
rect 8527 10217 8539 10251
rect 8481 10211 8539 10217
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 9640 10220 10425 10248
rect 9640 10208 9646 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 10413 10211 10471 10217
rect 12912 10220 13829 10248
rect 5350 10180 5356 10192
rect 5263 10152 5356 10180
rect 5350 10140 5356 10152
rect 5408 10180 5414 10192
rect 5408 10152 6408 10180
rect 5408 10140 5414 10152
rect 6380 10124 6408 10152
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2038 10112 2044 10124
rect 1995 10084 2044 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10112 2746 10124
rect 3970 10112 3976 10124
rect 2740 10084 3976 10112
rect 2740 10072 2746 10084
rect 3970 10072 3976 10084
rect 4028 10112 4034 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 4028 10084 4261 10112
rect 4028 10072 4034 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4706 10112 4712 10124
rect 4667 10084 4712 10112
rect 4249 10075 4307 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5684 10084 6285 10112
rect 5684 10072 5690 10084
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6822 10112 6828 10124
rect 6420 10084 6465 10112
rect 6783 10084 6828 10112
rect 6420 10072 6426 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7006 10112 7012 10124
rect 6967 10084 7012 10112
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 8260 10084 8309 10112
rect 8260 10072 8266 10084
rect 8297 10081 8309 10084
rect 8343 10112 8355 10115
rect 9858 10112 9864 10124
rect 8343 10084 9864 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10226 10112 10232 10124
rect 10187 10084 10232 10112
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12912 10121 12940 10220
rect 13817 10217 13829 10220
rect 13863 10248 13875 10251
rect 14734 10248 14740 10260
rect 13863 10220 14740 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 18414 10248 18420 10260
rect 17635 10220 18420 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 18564 10220 21281 10248
rect 18564 10208 18570 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 21269 10211 21327 10217
rect 21358 10208 21364 10260
rect 21416 10248 21422 10260
rect 21545 10251 21603 10257
rect 21545 10248 21557 10251
rect 21416 10220 21557 10248
rect 21416 10208 21422 10220
rect 21545 10217 21557 10220
rect 21591 10217 21603 10251
rect 22002 10248 22008 10260
rect 21963 10220 22008 10248
rect 21545 10211 21603 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 23014 10248 23020 10260
rect 22975 10220 23020 10248
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 17037 10183 17095 10189
rect 17037 10149 17049 10183
rect 17083 10180 17095 10183
rect 18524 10180 18552 10208
rect 17083 10152 18552 10180
rect 17083 10149 17095 10152
rect 17037 10143 17095 10149
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12400 10084 12909 10112
rect 12400 10072 12406 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 15562 10112 15568 10124
rect 15523 10084 15568 10112
rect 13081 10075 13139 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12986 10044 12992 10056
rect 12207 10016 12992 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 1872 9976 1900 10007
rect 12986 10004 12992 10016
rect 13044 10044 13050 10056
rect 13096 10044 13124 10075
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 16850 10112 16856 10124
rect 16715 10084 16856 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 16850 10072 16856 10084
rect 16908 10112 16914 10124
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 16908 10084 17969 10112
rect 16908 10072 16914 10084
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 18322 10112 18328 10124
rect 18283 10084 18328 10112
rect 17957 10075 18015 10081
rect 18322 10072 18328 10084
rect 18380 10112 18386 10124
rect 18785 10115 18843 10121
rect 18785 10112 18797 10115
rect 18380 10084 18797 10112
rect 18380 10072 18386 10084
rect 18785 10081 18797 10084
rect 18831 10081 18843 10115
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 18785 10075 18843 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 22646 10112 22652 10124
rect 22607 10084 22652 10112
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 13044 10016 13124 10044
rect 13044 10004 13050 10016
rect 15010 10004 15016 10056
rect 15068 10044 15074 10056
rect 15286 10044 15292 10056
rect 15068 10016 15292 10044
rect 15068 10004 15074 10016
rect 15286 10004 15292 10016
rect 15344 10044 15350 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 15344 10016 15485 10044
rect 15344 10004 15350 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17460 10016 17785 10044
rect 17460 10004 17466 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 2866 9976 2872 9988
rect 1872 9948 2872 9976
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 7650 9936 7656 9988
rect 7708 9976 7714 9988
rect 8757 9979 8815 9985
rect 8757 9976 8769 9979
rect 7708 9948 8769 9976
rect 7708 9936 7714 9948
rect 8757 9945 8769 9948
rect 8803 9945 8815 9979
rect 8757 9939 8815 9945
rect 12529 9979 12587 9985
rect 12529 9945 12541 9979
rect 12575 9976 12587 9979
rect 12802 9976 12808 9988
rect 12575 9948 12808 9976
rect 12575 9945 12587 9948
rect 12529 9939 12587 9945
rect 12802 9936 12808 9948
rect 12860 9976 12866 9988
rect 13354 9976 13360 9988
rect 12860 9948 13360 9976
rect 12860 9936 12866 9948
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 17788 9976 17816 10007
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 17920 10016 18245 10044
rect 17920 10004 17926 10016
rect 18233 10013 18245 10016
rect 18279 10044 18291 10047
rect 19150 10044 19156 10056
rect 18279 10016 19156 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 19426 9976 19432 9988
rect 17788 9948 19432 9976
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 2958 9908 2964 9920
rect 2919 9880 2964 9908
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 7524 9880 7757 9908
rect 7524 9868 7530 9880
rect 7745 9877 7757 9880
rect 7791 9877 7803 9911
rect 9950 9908 9956 9920
rect 9911 9880 9956 9908
rect 7745 9871 7803 9877
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12952 9880 13185 9908
rect 12952 9868 12958 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 14826 9908 14832 9920
rect 14739 9880 14832 9908
rect 13173 9871 13231 9877
rect 14826 9868 14832 9880
rect 14884 9908 14890 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14884 9880 14933 9908
rect 14884 9868 14890 9880
rect 14921 9877 14933 9880
rect 14967 9908 14979 9911
rect 15286 9908 15292 9920
rect 14967 9880 15292 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15746 9908 15752 9920
rect 15707 9880 15752 9908
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 1104 9818 24656 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 24656 9818
rect 1104 9744 24656 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2682 9704 2688 9716
rect 2087 9676 2688 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8481 9707 8539 9713
rect 8481 9704 8493 9707
rect 8260 9676 8493 9704
rect 8260 9664 8266 9676
rect 8481 9673 8493 9676
rect 8527 9673 8539 9707
rect 8481 9667 8539 9673
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 16850 9704 16856 9716
rect 15068 9676 16856 9704
rect 15068 9664 15074 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 17402 9704 17408 9716
rect 17363 9676 17408 9704
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 18601 9707 18659 9713
rect 18601 9704 18613 9707
rect 18472 9676 18613 9704
rect 18472 9664 18478 9676
rect 18601 9673 18613 9676
rect 18647 9673 18659 9707
rect 18601 9667 18659 9673
rect 20349 9707 20407 9713
rect 20349 9673 20361 9707
rect 20395 9704 20407 9707
rect 20530 9704 20536 9716
rect 20395 9676 20536 9704
rect 20395 9673 20407 9676
rect 20349 9667 20407 9673
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 22465 9707 22523 9713
rect 22465 9704 22477 9707
rect 20680 9676 22477 9704
rect 20680 9664 20686 9676
rect 22465 9673 22477 9676
rect 22511 9673 22523 9707
rect 22465 9667 22523 9673
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 23382 9704 23388 9716
rect 22704 9676 23388 9704
rect 22704 9664 22710 9676
rect 23382 9664 23388 9676
rect 23440 9704 23446 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23440 9676 23857 9704
rect 23440 9664 23446 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 6089 9639 6147 9645
rect 6089 9605 6101 9639
rect 6135 9636 6147 9639
rect 18325 9639 18383 9645
rect 6135 9608 7144 9636
rect 6135 9605 6147 9608
rect 6089 9599 6147 9605
rect 7116 9580 7144 9608
rect 18325 9605 18337 9639
rect 18371 9636 18383 9639
rect 18506 9636 18512 9648
rect 18371 9608 18512 9636
rect 18371 9605 18383 9608
rect 18325 9599 18383 9605
rect 18506 9596 18512 9608
rect 18564 9596 18570 9648
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2958 9568 2964 9580
rect 2455 9540 2964 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 5684 9540 7021 9568
rect 5684 9528 5690 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7156 9540 7941 9568
rect 7156 9528 7162 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12250 9568 12256 9580
rect 12115 9540 12256 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12250 9528 12256 9540
rect 12308 9568 12314 9580
rect 12894 9568 12900 9580
rect 12308 9540 12900 9568
rect 12308 9528 12314 9540
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 14936 9540 15424 9568
rect 14936 9512 14964 9540
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9500 6515 9503
rect 7466 9500 7472 9512
rect 6503 9472 7472 9500
rect 6503 9469 6515 9472
rect 6457 9463 6515 9469
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 1854 9364 1860 9376
rect 1719 9336 1860 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2700 9364 2728 9463
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 10134 9500 10140 9512
rect 10095 9472 10140 9500
rect 8021 9463 8079 9469
rect 3970 9392 3976 9444
rect 4028 9392 4034 9444
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 8036 9432 8064 9463
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 10502 9500 10508 9512
rect 10192 9472 10508 9500
rect 10192 9460 10198 9472
rect 10502 9460 10508 9472
rect 10560 9500 10566 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10560 9472 10885 9500
rect 10560 9460 10566 9472
rect 10873 9469 10885 9472
rect 10919 9500 10931 9503
rect 11241 9503 11299 9509
rect 11241 9500 11253 9503
rect 10919 9472 11253 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 11241 9469 11253 9472
rect 11287 9469 11299 9503
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 11241 9463 11299 9469
rect 11624 9472 12633 9500
rect 9490 9432 9496 9444
rect 6880 9404 8064 9432
rect 9451 9404 9496 9432
rect 6880 9392 6886 9404
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 10318 9392 10324 9444
rect 10376 9432 10382 9444
rect 11624 9441 11652 9472
rect 12621 9469 12633 9472
rect 12667 9469 12679 9503
rect 14918 9500 14924 9512
rect 14879 9472 14924 9500
rect 12621 9463 12679 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15286 9500 15292 9512
rect 15247 9472 15292 9500
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15396 9509 15424 9540
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 16666 9500 16672 9512
rect 16627 9472 16672 9500
rect 15381 9463 15439 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 20162 9500 20168 9512
rect 20123 9472 20168 9500
rect 20162 9460 20168 9472
rect 20220 9500 20226 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20220 9472 20637 9500
rect 20220 9460 20226 9472
rect 20625 9469 20637 9472
rect 20671 9500 20683 9503
rect 21266 9500 21272 9512
rect 20671 9472 21272 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 22189 9503 22247 9509
rect 22189 9500 22201 9503
rect 21836 9472 22201 9500
rect 11609 9435 11667 9441
rect 11609 9432 11621 9435
rect 10376 9404 11621 9432
rect 10376 9392 10382 9404
rect 11609 9401 11621 9404
rect 11655 9401 11667 9435
rect 11609 9395 11667 9401
rect 13354 9392 13360 9444
rect 13412 9392 13418 9444
rect 14642 9432 14648 9444
rect 14603 9404 14648 9432
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 15838 9432 15844 9444
rect 15799 9404 15844 9432
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 18230 9392 18236 9444
rect 18288 9432 18294 9444
rect 19061 9435 19119 9441
rect 19061 9432 19073 9435
rect 18288 9404 19073 9432
rect 18288 9392 18294 9404
rect 19061 9401 19073 9404
rect 19107 9432 19119 9435
rect 21174 9432 21180 9444
rect 19107 9404 21180 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 21836 9376 21864 9472
rect 22189 9469 22201 9472
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9469 22339 9503
rect 22281 9463 22339 9469
rect 3694 9364 3700 9376
rect 2700 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 5902 9364 5908 9376
rect 5767 9336 5908 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 9217 9367 9275 9373
rect 9217 9333 9229 9367
rect 9263 9364 9275 9367
rect 9674 9364 9680 9376
rect 9263 9336 9680 9364
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10284 9336 10609 9364
rect 10284 9324 10290 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 11054 9364 11060 9376
rect 10643 9336 11060 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15562 9364 15568 9376
rect 15252 9336 15568 9364
rect 15252 9324 15258 9336
rect 15562 9324 15568 9336
rect 15620 9364 15626 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 15620 9336 16129 9364
rect 15620 9324 15626 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 21082 9364 21088 9376
rect 21043 9336 21088 9364
rect 16117 9327 16175 9333
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 21818 9364 21824 9376
rect 21779 9336 21824 9364
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 22296 9364 22324 9463
rect 23106 9364 23112 9376
rect 22296 9336 23112 9364
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 1104 9274 24656 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 24656 9274
rect 1104 9200 24656 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3421 9163 3479 9169
rect 3421 9160 3433 9163
rect 2924 9132 3433 9160
rect 2924 9120 2930 9132
rect 3421 9129 3433 9132
rect 3467 9129 3479 9163
rect 3421 9123 3479 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4120 9132 4261 9160
rect 4120 9120 4126 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5684 9132 5825 9160
rect 5684 9120 5690 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5960 9132 6193 9160
rect 5960 9120 5966 9132
rect 6181 9129 6193 9132
rect 6227 9160 6239 9163
rect 6822 9160 6828 9172
rect 6227 9132 6828 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 6822 9120 6828 9132
rect 6880 9160 6886 9172
rect 9309 9163 9367 9169
rect 6880 9132 6960 9160
rect 6880 9120 6886 9132
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 4614 9092 4620 9104
rect 3191 9064 4620 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 6932 9101 6960 9132
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9490 9160 9496 9172
rect 9355 9132 9496 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15010 9160 15016 9172
rect 14967 9132 15016 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 17773 9163 17831 9169
rect 17773 9129 17785 9163
rect 17819 9160 17831 9163
rect 18322 9160 18328 9172
rect 17819 9132 18328 9160
rect 17819 9129 17831 9132
rect 17773 9123 17831 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 6917 9095 6975 9101
rect 6917 9061 6929 9095
rect 6963 9061 6975 9095
rect 9508 9092 9536 9120
rect 10410 9092 10416 9104
rect 9508 9064 10416 9092
rect 6917 9055 6975 9061
rect 10410 9052 10416 9064
rect 10468 9092 10474 9104
rect 17405 9095 17463 9101
rect 10468 9064 10916 9092
rect 10468 9052 10474 9064
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 5074 9024 5080 9036
rect 5035 8996 5080 9024
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 5960 8996 7021 9024
rect 5960 8984 5966 8996
rect 7009 8993 7021 8996
rect 7055 9024 7067 9027
rect 7650 9024 7656 9036
rect 7055 8996 7656 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 8260 8996 8585 9024
rect 8260 8984 8266 8996
rect 8573 8993 8585 8996
rect 8619 8993 8631 9027
rect 10502 9024 10508 9036
rect 10463 8996 10508 9024
rect 8573 8987 8631 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10888 9033 10916 9064
rect 17405 9061 17417 9095
rect 17451 9092 17463 9095
rect 17862 9092 17868 9104
rect 17451 9064 17868 9092
rect 17451 9061 17463 9064
rect 17405 9055 17463 9061
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 22278 9052 22284 9104
rect 22336 9052 22342 9104
rect 23382 9052 23388 9104
rect 23440 9092 23446 9104
rect 23477 9095 23535 9101
rect 23477 9092 23489 9095
rect 23440 9064 23489 9092
rect 23440 9052 23446 9064
rect 23477 9061 23489 9064
rect 23523 9061 23535 9095
rect 23477 9055 23535 9061
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 10919 8996 11345 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 12250 9024 12256 9036
rect 12211 8996 12256 9024
rect 11333 8987 11391 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 9024 13050 9036
rect 14642 9024 14648 9036
rect 13044 8996 14648 9024
rect 13044 8984 13050 8996
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 15562 9024 15568 9036
rect 15523 8996 15568 9024
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 18196 8996 18613 9024
rect 18196 8984 18202 8996
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 10318 8956 10324 8968
rect 3752 8928 4154 8956
rect 10279 8928 10324 8956
rect 3752 8916 3758 8928
rect 2777 8891 2835 8897
rect 2777 8857 2789 8891
rect 2823 8888 2835 8891
rect 3970 8888 3976 8900
rect 2823 8860 3976 8888
rect 2823 8857 2835 8860
rect 2777 8851 2835 8857
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 4126 8888 4154 8928
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 10778 8956 10784 8968
rect 10739 8928 10784 8956
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 12400 8928 13277 8956
rect 12400 8916 12406 8928
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 14148 8928 15485 8956
rect 14148 8916 14154 8928
rect 15473 8925 15485 8928
rect 15519 8956 15531 8959
rect 16666 8956 16672 8968
rect 15519 8928 16672 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21232 8928 21465 8956
rect 21232 8916 21238 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21726 8956 21732 8968
rect 21687 8928 21732 8956
rect 21453 8919 21511 8925
rect 4709 8891 4767 8897
rect 4709 8888 4721 8891
rect 4126 8860 4721 8888
rect 4709 8857 4721 8860
rect 4755 8888 4767 8891
rect 6641 8891 6699 8897
rect 4755 8860 6592 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 1854 8820 1860 8832
rect 1815 8792 1860 8820
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 5224 8792 5273 8820
rect 5224 8780 5230 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 6564 8820 6592 8860
rect 6641 8857 6653 8891
rect 6687 8888 6699 8891
rect 7006 8888 7012 8900
rect 6687 8860 7012 8888
rect 6687 8857 6699 8860
rect 6641 8851 6699 8857
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 12529 8891 12587 8897
rect 12529 8888 12541 8891
rect 11940 8860 12541 8888
rect 11940 8848 11946 8860
rect 12529 8857 12541 8860
rect 12575 8857 12587 8891
rect 12529 8851 12587 8857
rect 18233 8891 18291 8897
rect 18233 8857 18245 8891
rect 18279 8888 18291 8891
rect 19242 8888 19248 8900
rect 18279 8860 19248 8888
rect 18279 8857 18291 8860
rect 18233 8851 18291 8857
rect 19242 8848 19248 8860
rect 19300 8848 19306 8900
rect 6914 8820 6920 8832
rect 6564 8792 6920 8820
rect 5261 8783 5319 8789
rect 6914 8780 6920 8792
rect 6972 8820 6978 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 6972 8792 7941 8820
rect 6972 8780 6978 8792
rect 7929 8789 7941 8792
rect 7975 8820 7987 8823
rect 8662 8820 8668 8832
rect 7975 8792 8668 8820
rect 7975 8789 7987 8792
rect 7929 8783 7987 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 10594 8820 10600 8832
rect 8803 8792 10600 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 19484 8792 19533 8820
rect 19484 8780 19490 8792
rect 19521 8789 19533 8792
rect 19567 8789 19579 8823
rect 21468 8820 21496 8919
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 22738 8820 22744 8832
rect 21468 8792 22744 8820
rect 19521 8783 19579 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 1104 8730 24656 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 24656 8730
rect 1104 8656 24656 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2041 8619 2099 8625
rect 2041 8616 2053 8619
rect 1728 8588 2053 8616
rect 1728 8576 1734 8588
rect 2041 8585 2053 8588
rect 2087 8585 2099 8619
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 2041 8579 2099 8585
rect 3510 8576 3516 8588
rect 3568 8616 3574 8628
rect 4046 8619 4104 8625
rect 4046 8616 4058 8619
rect 3568 8588 4058 8616
rect 3568 8576 3574 8588
rect 4046 8585 4058 8588
rect 4092 8585 4104 8619
rect 4046 8579 4104 8585
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 10318 8616 10324 8628
rect 9447 8588 10324 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 10744 8588 12817 8616
rect 10744 8576 10750 8588
rect 12805 8585 12817 8588
rect 12851 8585 12863 8619
rect 12805 8579 12863 8585
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12952 8588 13093 8616
rect 12952 8576 12958 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16666 8616 16672 8628
rect 16439 8588 16672 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 20809 8619 20867 8625
rect 20809 8616 20821 8619
rect 16908 8588 20821 8616
rect 16908 8576 16914 8588
rect 20809 8585 20821 8588
rect 20855 8585 20867 8619
rect 20809 8579 20867 8585
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3191 8452 5212 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 5184 8424 5212 8452
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6972 8452 7021 8480
rect 6972 8440 6978 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 7708 8452 9045 8480
rect 7708 8440 7714 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 15470 8480 15476 8492
rect 15431 8452 15476 8480
rect 9033 8443 9091 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 18138 8440 18144 8492
rect 18196 8480 18202 8492
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 18196 8452 20269 8480
rect 18196 8440 18202 8452
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 20824 8480 20852 8579
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 21140 8588 21833 8616
rect 21140 8576 21146 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 21545 8483 21603 8489
rect 21545 8480 21557 8483
rect 20824 8452 21557 8480
rect 20257 8443 20315 8449
rect 21545 8449 21557 8452
rect 21591 8480 21603 8483
rect 21818 8480 21824 8492
rect 21591 8452 21824 8480
rect 21591 8449 21603 8452
rect 21545 8443 21603 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 1854 8412 1860 8424
rect 1627 8384 1860 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3752 8384 3801 8412
rect 3752 8372 3758 8384
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 5166 8372 5172 8424
rect 5224 8372 5230 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 6822 8412 6828 8424
rect 5859 8384 6828 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 9674 8412 9680 8424
rect 9635 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9858 8412 9864 8424
rect 9819 8384 9864 8412
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10410 8372 10416 8424
rect 10468 8412 10474 8424
rect 10597 8415 10655 8421
rect 10468 8384 10513 8412
rect 10468 8372 10474 8384
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10778 8412 10784 8424
rect 10643 8384 10784 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10778 8372 10784 8384
rect 10836 8412 10842 8424
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 10836 8384 11376 8412
rect 10836 8372 10842 8384
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 7282 8344 7288 8356
rect 6503 8316 7288 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 7926 8304 7932 8356
rect 7984 8304 7990 8356
rect 11348 8288 11376 8384
rect 11992 8384 12633 8412
rect 1670 8236 1676 8288
rect 1728 8276 1734 8288
rect 1765 8279 1823 8285
rect 1765 8276 1777 8279
rect 1728 8248 1777 8276
rect 1728 8236 1734 8248
rect 1765 8245 1777 8248
rect 1811 8245 1823 8279
rect 1765 8239 1823 8245
rect 2501 8279 2559 8285
rect 2501 8245 2513 8279
rect 2547 8276 2559 8279
rect 2958 8276 2964 8288
rect 2547 8248 2964 8276
rect 2547 8245 2559 8248
rect 2501 8239 2559 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 10192 8248 10885 8276
rect 10192 8236 10198 8248
rect 10873 8245 10885 8248
rect 10919 8245 10931 8279
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 10873 8239 10931 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11992 8285 12020 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 12621 8375 12679 8381
rect 14016 8384 14381 8412
rect 14016 8288 14044 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 15838 8412 15844 8424
rect 15799 8384 15844 8412
rect 14369 8375 14427 8381
rect 15838 8372 15844 8384
rect 15896 8412 15902 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 15896 8384 16681 8412
rect 15896 8372 15902 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 18230 8412 18236 8424
rect 18191 8384 18236 8412
rect 16669 8375 16727 8381
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 21637 8415 21695 8421
rect 21637 8381 21649 8415
rect 21683 8412 21695 8415
rect 21683 8384 22508 8412
rect 21683 8381 21695 8384
rect 21637 8375 21695 8381
rect 17221 8347 17279 8353
rect 17221 8344 17233 8347
rect 16040 8316 17233 8344
rect 16040 8288 16068 8316
rect 17221 8313 17233 8316
rect 17267 8313 17279 8347
rect 17221 8307 17279 8313
rect 17681 8347 17739 8353
rect 17681 8313 17693 8347
rect 17727 8344 17739 8347
rect 18506 8344 18512 8356
rect 17727 8316 18512 8344
rect 17727 8313 17739 8316
rect 17681 8307 17739 8313
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 19242 8304 19248 8356
rect 19300 8304 19306 8356
rect 22480 8353 22508 8384
rect 22465 8347 22523 8353
rect 22465 8313 22477 8347
rect 22511 8344 22523 8347
rect 24486 8344 24492 8356
rect 22511 8316 24492 8344
rect 22511 8313 22523 8316
rect 22465 8307 22523 8313
rect 24486 8304 24492 8316
rect 24544 8304 24550 8356
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11756 8248 11989 8276
rect 11756 8236 11762 8248
rect 11977 8245 11989 8248
rect 12023 8245 12035 8279
rect 13998 8276 14004 8288
rect 13959 8248 14004 8276
rect 11977 8239 12035 8245
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 14737 8279 14795 8285
rect 14737 8245 14749 8279
rect 14783 8276 14795 8279
rect 14826 8276 14832 8288
rect 14783 8248 14832 8276
rect 14783 8245 14795 8248
rect 14737 8239 14795 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 16022 8276 16028 8288
rect 15983 8248 16028 8276
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 21269 8279 21327 8285
rect 21269 8245 21281 8279
rect 21315 8276 21327 8279
rect 21726 8276 21732 8288
rect 21315 8248 21732 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 22738 8276 22744 8288
rect 22699 8248 22744 8276
rect 22738 8236 22744 8248
rect 22796 8236 22802 8288
rect 1104 8186 24656 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 24656 8186
rect 1104 8112 24656 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3694 8072 3700 8084
rect 3467 8044 3700 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4028 8044 4445 8072
rect 4028 8032 4034 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 5074 8072 5080 8084
rect 5035 8044 5080 8072
rect 4433 8035 4491 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7926 8072 7932 8084
rect 7331 8044 7932 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 10778 8072 10784 8084
rect 9355 8044 10784 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 12342 8072 12348 8084
rect 12303 8044 12348 8072
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12986 8072 12992 8084
rect 12759 8044 12992 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 19300 8044 21281 8072
rect 19300 8032 19306 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 21637 8075 21695 8081
rect 21637 8041 21649 8075
rect 21683 8072 21695 8075
rect 22278 8072 22284 8084
rect 21683 8044 22284 8072
rect 21683 8041 21695 8044
rect 21637 8035 21695 8041
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 22370 8032 22376 8084
rect 22428 8072 22434 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 22428 8044 22569 8072
rect 22428 8032 22434 8044
rect 22557 8041 22569 8044
rect 22603 8041 22615 8075
rect 22557 8035 22615 8041
rect 5092 8004 5120 8032
rect 7466 8004 7472 8016
rect 5092 7976 7472 8004
rect 7466 7964 7472 7976
rect 7524 8004 7530 8016
rect 8297 8007 8355 8013
rect 7524 7976 7788 8004
rect 7524 7964 7530 7976
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 4120 7908 4261 7936
rect 4120 7896 4126 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 6822 7936 6828 7948
rect 6783 7908 6828 7936
rect 4249 7899 4307 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7760 7945 7788 7976
rect 8297 7973 8309 8007
rect 8343 8004 8355 8007
rect 8754 8004 8760 8016
rect 8343 7976 8760 8004
rect 8343 7973 8355 7976
rect 8297 7967 8355 7973
rect 8754 7964 8760 7976
rect 8812 8004 8818 8016
rect 9858 8004 9864 8016
rect 8812 7976 9864 8004
rect 8812 7964 8818 7976
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10134 8004 10140 8016
rect 10095 7976 10140 8004
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10594 7964 10600 8016
rect 10652 7964 10658 8016
rect 16209 8007 16267 8013
rect 16209 7973 16221 8007
rect 16255 8004 16267 8007
rect 16255 7976 17448 8004
rect 16255 7973 16267 7976
rect 16209 7967 16267 7973
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7936 7803 7939
rect 8202 7936 8208 7948
rect 7791 7908 8208 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 8202 7896 8208 7908
rect 8260 7936 8266 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8260 7908 8585 7936
rect 8260 7896 8266 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 14967 7908 15485 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 15473 7905 15485 7908
rect 15519 7936 15531 7939
rect 15746 7936 15752 7948
rect 15519 7908 15752 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 16080 7908 16589 7936
rect 16080 7896 16086 7908
rect 16577 7905 16589 7908
rect 16623 7936 16635 7939
rect 16942 7936 16948 7948
rect 16623 7908 16948 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 17420 7945 17448 7976
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7936 17463 7939
rect 17451 7908 18092 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 8720 7840 9873 7868
rect 8720 7828 8726 7840
rect 9861 7837 9873 7840
rect 9907 7868 9919 7871
rect 10226 7868 10232 7880
rect 9907 7840 10232 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 10560 7840 11897 7868
rect 10560 7828 10566 7840
rect 11885 7837 11897 7840
rect 11931 7837 11943 7871
rect 11885 7831 11943 7837
rect 18064 7800 18092 7908
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 19337 7939 19395 7945
rect 19337 7936 19349 7939
rect 18380 7908 19349 7936
rect 18380 7896 18386 7908
rect 19337 7905 19349 7908
rect 19383 7936 19395 7939
rect 19426 7936 19432 7948
rect 19383 7908 19432 7936
rect 19383 7905 19395 7908
rect 19337 7899 19395 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 20438 7896 20444 7948
rect 20496 7936 20502 7948
rect 21085 7939 21143 7945
rect 21085 7936 21097 7939
rect 20496 7908 21097 7936
rect 20496 7896 20502 7908
rect 21085 7905 21097 7908
rect 21131 7936 21143 7939
rect 22097 7939 22155 7945
rect 22097 7936 22109 7939
rect 21131 7908 22109 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 22097 7905 22109 7908
rect 22143 7936 22155 7939
rect 22388 7936 22416 8032
rect 23109 7939 23167 7945
rect 23109 7936 23121 7939
rect 22143 7908 23121 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 23109 7905 23121 7908
rect 23155 7936 23167 7939
rect 23198 7936 23204 7948
rect 23155 7908 23204 7936
rect 23155 7905 23167 7908
rect 23109 7899 23167 7905
rect 23198 7896 23204 7908
rect 23256 7896 23262 7948
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18690 7868 18696 7880
rect 18463 7840 18696 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19024 7840 19257 7868
rect 19024 7828 19030 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 18598 7800 18604 7812
rect 18064 7772 18604 7800
rect 18598 7760 18604 7772
rect 18656 7800 18662 7812
rect 20257 7803 20315 7809
rect 20257 7800 20269 7803
rect 18656 7772 20269 7800
rect 18656 7760 18662 7772
rect 20257 7769 20269 7772
rect 20303 7769 20315 7803
rect 20257 7763 20315 7769
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 2222 7732 2228 7744
rect 2087 7704 2228 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2222 7692 2228 7704
rect 2280 7732 2286 7744
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2280 7704 2605 7732
rect 2280 7692 2286 7704
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 2593 7695 2651 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 14090 7732 14096 7744
rect 14051 7704 14096 7732
rect 14090 7692 14096 7704
rect 14148 7732 14154 7744
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 14148 7704 15669 7732
rect 14148 7692 14154 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18196 7704 18705 7732
rect 18196 7692 18202 7704
rect 18693 7701 18705 7704
rect 18739 7701 18751 7735
rect 23290 7732 23296 7744
rect 23251 7704 23296 7732
rect 18693 7695 18751 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 1104 7642 24656 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 24656 7642
rect 1104 7568 24656 7590
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 23198 7528 23204 7540
rect 23159 7500 23204 7528
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 7193 7463 7251 7469
rect 7193 7429 7205 7463
rect 7239 7460 7251 7463
rect 7239 7432 9444 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2280 7364 2881 7392
rect 2280 7352 2286 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2406 7324 2412 7336
rect 1719 7296 2412 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4062 7324 4068 7336
rect 3975 7296 4068 7324
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 6273 7327 6331 7333
rect 4120 7296 4660 7324
rect 4120 7284 4126 7296
rect 1946 7256 1952 7268
rect 1907 7228 1952 7256
rect 1946 7216 1952 7228
rect 2004 7216 2010 7268
rect 2424 7256 2452 7284
rect 2424 7228 3556 7256
rect 3528 7197 3556 7228
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 3694 7188 3700 7200
rect 3559 7160 3700 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4632 7197 4660 7296
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 6822 7324 6828 7336
rect 6319 7296 6828 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 6822 7284 6828 7296
rect 6880 7324 6886 7336
rect 7650 7324 7656 7336
rect 6880 7296 7656 7324
rect 6880 7284 6886 7296
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 8754 7324 8760 7336
rect 8715 7296 8760 7324
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9416 7324 9444 7432
rect 18506 7420 18512 7472
rect 18564 7460 18570 7472
rect 19337 7463 19395 7469
rect 19337 7460 19349 7463
rect 18564 7432 19349 7460
rect 18564 7420 18570 7432
rect 19337 7429 19349 7432
rect 19383 7429 19395 7463
rect 19337 7423 19395 7429
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 14090 7392 14096 7404
rect 14051 7364 14096 7392
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 16298 7392 16304 7404
rect 15488 7364 16304 7392
rect 9674 7324 9680 7336
rect 9263 7296 9680 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9674 7284 9680 7296
rect 9732 7324 9738 7336
rect 10134 7324 10140 7336
rect 9732 7296 10140 7324
rect 9732 7284 9738 7296
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10376 7296 10701 7324
rect 10376 7284 10382 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 14274 7324 14280 7336
rect 10689 7287 10747 7293
rect 13372 7296 14280 7324
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7340 7228 8892 7256
rect 7340 7216 7346 7228
rect 4249 7191 4307 7197
rect 4249 7188 4261 7191
rect 3844 7160 4261 7188
rect 3844 7148 3850 7160
rect 4249 7157 4261 7160
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7188 4675 7191
rect 4982 7188 4988 7200
rect 4663 7160 4988 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13372 7197 13400 7296
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 13817 7259 13875 7265
rect 13817 7225 13829 7259
rect 13863 7256 13875 7259
rect 14752 7256 14780 7287
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 14884 7296 14929 7324
rect 14884 7284 14890 7296
rect 15488 7256 15516 7364
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 17000 7364 18245 7392
rect 17000 7352 17006 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 13863 7228 15516 7256
rect 15948 7296 16405 7324
rect 13863 7225 13875 7228
rect 13817 7219 13875 7225
rect 15948 7200 15976 7296
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18598 7324 18604 7336
rect 18463 7296 18604 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 18782 7284 18788 7336
rect 18840 7324 18846 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18840 7296 18889 7324
rect 18840 7284 18846 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 20073 7327 20131 7333
rect 19024 7296 19069 7324
rect 19024 7284 19030 7296
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 20806 7324 20812 7336
rect 20119 7296 20812 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 21542 7324 21548 7336
rect 21503 7296 21548 7324
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 17310 7216 17316 7268
rect 17368 7256 17374 7268
rect 17681 7259 17739 7265
rect 17681 7256 17693 7259
rect 17368 7228 17693 7256
rect 17368 7216 17374 7228
rect 17681 7225 17693 7228
rect 17727 7256 17739 7259
rect 18800 7256 18828 7284
rect 17727 7228 18828 7256
rect 17727 7225 17739 7228
rect 17681 7219 17739 7225
rect 21726 7216 21732 7268
rect 21784 7216 21790 7268
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 13044 7160 13369 7188
rect 13044 7148 13050 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13357 7151 13415 7157
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 15068 7160 15301 7188
rect 15068 7148 15074 7160
rect 15289 7157 15301 7160
rect 15335 7157 15347 7191
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 15289 7151 15347 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 1104 7098 24656 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 24656 7098
rect 1104 7024 24656 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3602 6984 3608 6996
rect 2648 6956 3608 6984
rect 2648 6944 2654 6956
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10502 6984 10508 6996
rect 9999 6956 10508 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 14185 6987 14243 6993
rect 14185 6953 14197 6987
rect 14231 6984 14243 6987
rect 14826 6984 14832 6996
rect 14231 6956 14832 6984
rect 14231 6953 14243 6956
rect 14185 6947 14243 6953
rect 14826 6944 14832 6956
rect 14884 6984 14890 6996
rect 16942 6984 16948 6996
rect 14884 6956 16528 6984
rect 16903 6956 16948 6984
rect 14884 6944 14890 6956
rect 2958 6916 2964 6928
rect 2332 6888 2964 6916
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 1946 6848 1952 6860
rect 1811 6820 1952 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 2332 6857 2360 6888
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 5350 6916 5356 6928
rect 4571 6888 5356 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 5350 6876 5356 6888
rect 5408 6916 5414 6928
rect 5408 6888 5488 6916
rect 5408 6876 5414 6888
rect 5460 6857 5488 6888
rect 5810 6876 5816 6928
rect 5868 6876 5874 6928
rect 10226 6916 10232 6928
rect 10187 6888 10232 6916
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 10318 6876 10324 6928
rect 10376 6916 10382 6928
rect 10597 6919 10655 6925
rect 10597 6916 10609 6919
rect 10376 6888 10609 6916
rect 10376 6876 10382 6888
rect 10597 6885 10609 6888
rect 10643 6885 10655 6919
rect 11882 6916 11888 6928
rect 11843 6888 11888 6916
rect 10597 6879 10655 6885
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 12342 6876 12348 6928
rect 12400 6876 12406 6928
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 15473 6919 15531 6925
rect 15473 6916 15485 6919
rect 14332 6888 15485 6916
rect 14332 6876 14338 6888
rect 15473 6885 15485 6888
rect 15519 6885 15531 6919
rect 15473 6879 15531 6885
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6914 6848 6920 6860
rect 6227 6820 6920 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7926 6848 7932 6860
rect 7887 6820 7932 6848
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 10244 6848 10272 6876
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 10244 6820 11621 6848
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 13998 6848 14004 6860
rect 13679 6820 14004 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 11624 6780 11652 6811
rect 13998 6808 14004 6820
rect 14056 6848 14062 6860
rect 16500 6857 16528 6956
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17957 6987 18015 6993
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18598 6984 18604 6996
rect 18003 6956 18604 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 17405 6919 17463 6925
rect 17405 6885 17417 6919
rect 17451 6916 17463 6919
rect 17770 6916 17776 6928
rect 17451 6888 17776 6916
rect 17451 6885 17463 6888
rect 17405 6879 17463 6885
rect 17770 6876 17776 6888
rect 17828 6916 17834 6928
rect 18966 6916 18972 6928
rect 17828 6888 18972 6916
rect 17828 6876 17834 6888
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14056 6820 14565 6848
rect 14056 6808 14062 6820
rect 14553 6817 14565 6820
rect 14599 6848 14611 6851
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 14599 6820 16129 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 18322 6848 18328 6860
rect 16724 6820 18328 6848
rect 16724 6808 16730 6820
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 18662 6857 18690 6888
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 20533 6919 20591 6925
rect 20533 6885 20545 6919
rect 20579 6916 20591 6919
rect 21542 6916 21548 6928
rect 20579 6888 21548 6916
rect 20579 6885 20591 6888
rect 20533 6879 20591 6885
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 18647 6851 18705 6857
rect 18647 6817 18659 6851
rect 18693 6817 18705 6851
rect 18782 6848 18788 6860
rect 18743 6820 18788 6848
rect 18647 6811 18705 6817
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 19886 6848 19892 6860
rect 19843 6820 19892 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 22922 6808 22928 6860
rect 22980 6808 22986 6860
rect 12618 6780 12624 6792
rect 11624 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 15930 6780 15936 6792
rect 15620 6752 15936 6780
rect 15620 6740 15626 6752
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16356 6752 16405 6780
rect 16356 6740 16362 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 18138 6780 18144 6792
rect 18099 6752 18144 6780
rect 16393 6743 16451 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 21082 6740 21088 6792
rect 21140 6780 21146 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 21140 6752 21557 6780
rect 21140 6740 21146 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21818 6780 21824 6792
rect 21779 6752 21824 6780
rect 21545 6743 21603 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 23566 6780 23572 6792
rect 23527 6752 23572 6780
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 1688 6644 1716 6740
rect 2682 6712 2688 6724
rect 2643 6684 2688 6712
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 1688 6616 3249 6644
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3237 6607 3295 6613
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7558 6644 7564 6656
rect 7147 6616 7564 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7558 6604 7564 6616
rect 7616 6644 7622 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7616 6616 7849 6644
rect 7616 6604 7622 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 19150 6644 19156 6656
rect 19111 6616 19156 6644
rect 7837 6607 7895 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6644 21327 6647
rect 22002 6644 22008 6656
rect 21315 6616 22008 6644
rect 21315 6613 21327 6616
rect 21269 6607 21327 6613
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 1104 6554 24656 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 24656 6554
rect 1104 6480 24656 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 3786 6440 3792 6452
rect 1811 6412 3792 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 6914 6440 6920 6452
rect 4939 6412 6920 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12618 6440 12624 6452
rect 12579 6412 12624 6440
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 17310 6440 17316 6452
rect 17271 6412 17316 6440
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 18138 6440 18144 6452
rect 17727 6412 18144 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 21085 6443 21143 6449
rect 21085 6409 21097 6443
rect 21131 6440 21143 6443
rect 21818 6440 21824 6452
rect 21131 6412 21824 6440
rect 21131 6409 21143 6412
rect 21085 6403 21143 6409
rect 21818 6400 21824 6412
rect 21876 6440 21882 6452
rect 22557 6443 22615 6449
rect 22557 6440 22569 6443
rect 21876 6412 22569 6440
rect 21876 6400 21882 6412
rect 22557 6409 22569 6412
rect 22603 6409 22615 6443
rect 22557 6403 22615 6409
rect 22922 6400 22928 6452
rect 22980 6440 22986 6452
rect 23109 6443 23167 6449
rect 23109 6440 23121 6443
rect 22980 6412 23121 6440
rect 22980 6400 22986 6412
rect 23109 6409 23121 6412
rect 23155 6440 23167 6443
rect 23290 6440 23296 6452
rect 23155 6412 23296 6440
rect 23155 6409 23167 6412
rect 23109 6403 23167 6409
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 11057 6375 11115 6381
rect 5859 6344 8892 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2682 6304 2688 6316
rect 2179 6276 2688 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 3752 6276 4445 6304
rect 3752 6264 3758 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 2406 6236 2412 6248
rect 2367 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 3786 6196 3792 6248
rect 3844 6196 3850 6248
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5040 6208 5273 6236
rect 5040 6196 5046 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5828 6236 5856 6335
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7616 6276 7941 6304
rect 7616 6264 7622 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 5307 6208 5856 6236
rect 7469 6239 7527 6245
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7650 6236 7656 6248
rect 7611 6208 7656 6236
rect 7469 6199 7527 6205
rect 5350 6128 5356 6180
rect 5408 6168 5414 6180
rect 7006 6168 7012 6180
rect 5408 6140 7012 6168
rect 5408 6128 5414 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 5040 6072 5457 6100
rect 5040 6060 5046 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 7484 6100 7512 6199
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 8018 6236 8024 6248
rect 7979 6208 8024 6236
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8864 6245 8892 6344
rect 11057 6341 11069 6375
rect 11103 6372 11115 6375
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 11103 6344 11529 6372
rect 11103 6341 11115 6344
rect 11057 6335 11115 6341
rect 11517 6341 11529 6344
rect 11563 6372 11575 6375
rect 12342 6372 12348 6384
rect 11563 6344 12348 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 15010 6304 15016 6316
rect 14507 6276 15016 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15562 6264 15568 6316
rect 15620 6304 15626 6316
rect 16761 6307 16819 6313
rect 16761 6304 16773 6307
rect 15620 6276 16773 6304
rect 15620 6264 15626 6276
rect 16761 6273 16773 6276
rect 16807 6273 16819 6307
rect 16761 6267 16819 6273
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18417 6307 18475 6313
rect 18417 6304 18429 6307
rect 18288 6276 18429 6304
rect 18288 6264 18294 6276
rect 18417 6273 18429 6276
rect 18463 6273 18475 6307
rect 18690 6304 18696 6316
rect 18651 6276 18696 6304
rect 18417 6267 18475 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 20806 6264 20812 6316
rect 20864 6304 20870 6316
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 20864 6276 21373 6304
rect 20864 6264 20870 6276
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8895 6208 9444 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 7926 6100 7932 6112
rect 6503 6072 7932 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 7926 6060 7932 6072
rect 7984 6100 7990 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 7984 6072 8585 6100
rect 7984 6060 7990 6072
rect 8573 6069 8585 6072
rect 8619 6100 8631 6103
rect 8754 6100 8760 6112
rect 8619 6072 8760 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9416 6109 9444 6208
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9824 6208 9965 6236
rect 9824 6196 9830 6208
rect 9953 6205 9965 6208
rect 9999 6236 10011 6239
rect 10410 6236 10416 6248
rect 9999 6208 10416 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 11790 6236 11796 6248
rect 11379 6208 11796 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8904 6072 9045 6100
rect 8904 6060 8910 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9447 6072 10149 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 10137 6069 10149 6072
rect 10183 6100 10195 6103
rect 11348 6100 11376 6199
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13786 6208 14105 6236
rect 10183 6072 11376 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 13786 6100 13814 6208
rect 14093 6205 14105 6208
rect 14139 6236 14151 6239
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 14139 6208 14749 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 21542 6236 21548 6248
rect 21503 6208 21548 6236
rect 14737 6199 14795 6205
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22281 6239 22339 6245
rect 22152 6208 22197 6236
rect 22152 6196 22158 6208
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 22830 6236 22836 6248
rect 22327 6208 22836 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 15470 6128 15476 6180
rect 15528 6128 15534 6180
rect 19150 6128 19156 6180
rect 19208 6128 19214 6180
rect 20438 6168 20444 6180
rect 20399 6140 20444 6168
rect 20438 6128 20444 6140
rect 20496 6128 20502 6180
rect 21082 6128 21088 6180
rect 21140 6168 21146 6180
rect 22738 6168 22744 6180
rect 21140 6140 22744 6168
rect 21140 6128 21146 6140
rect 22738 6128 22744 6140
rect 22796 6168 22802 6180
rect 23845 6171 23903 6177
rect 23845 6168 23857 6171
rect 22796 6140 23857 6168
rect 22796 6128 22802 6140
rect 23845 6137 23857 6140
rect 23891 6137 23903 6171
rect 23845 6131 23903 6137
rect 13688 6072 13814 6100
rect 13688 6060 13694 6072
rect 1104 6010 24656 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 24656 6010
rect 1104 5936 24656 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2222 5896 2228 5908
rect 1719 5868 2228 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2222 5856 2228 5868
rect 2280 5856 2286 5908
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 3050 5896 3056 5908
rect 2464 5868 3056 5896
rect 2464 5856 2470 5868
rect 3050 5856 3056 5868
rect 3108 5896 3114 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3108 5868 3433 5896
rect 3108 5856 3114 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 2958 5828 2964 5840
rect 2087 5800 2964 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 2958 5788 2964 5800
rect 3016 5828 3022 5840
rect 3145 5831 3203 5837
rect 3145 5828 3157 5831
rect 3016 5800 3157 5828
rect 3016 5788 3022 5800
rect 3145 5797 3157 5800
rect 3191 5797 3203 5831
rect 3145 5791 3203 5797
rect 2590 5760 2596 5772
rect 2551 5732 2596 5760
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 3436 5692 3464 5859
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 6638 5896 6644 5908
rect 3660 5868 6316 5896
rect 6599 5868 6644 5896
rect 3660 5856 3666 5868
rect 4982 5788 4988 5840
rect 5040 5788 5046 5840
rect 6288 5837 6316 5868
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 7708 5868 8585 5896
rect 7708 5856 7714 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 10134 5896 10140 5908
rect 10095 5868 10140 5896
rect 8573 5859 8631 5865
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 11790 5896 11796 5908
rect 11751 5868 11796 5896
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 15562 5896 15568 5908
rect 15523 5868 15568 5896
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 16298 5896 16304 5908
rect 15979 5868 16304 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 17770 5896 17776 5908
rect 17731 5868 17776 5896
rect 17770 5856 17776 5868
rect 17828 5856 17834 5908
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 18690 5896 18696 5908
rect 18555 5868 18696 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 18690 5856 18696 5868
rect 18748 5856 18754 5908
rect 19150 5856 19156 5908
rect 19208 5896 19214 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 19208 5868 19257 5896
rect 19208 5856 19214 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 20533 5899 20591 5905
rect 20533 5865 20545 5899
rect 20579 5896 20591 5899
rect 20806 5896 20812 5908
rect 20579 5868 20812 5896
rect 20579 5865 20591 5868
rect 20533 5859 20591 5865
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21600 5868 21925 5896
rect 21600 5856 21606 5868
rect 21913 5865 21925 5868
rect 21959 5896 21971 5899
rect 23109 5899 23167 5905
rect 23109 5896 23121 5899
rect 21959 5868 23121 5896
rect 21959 5865 21971 5868
rect 21913 5859 21971 5865
rect 23109 5865 23121 5868
rect 23155 5865 23167 5899
rect 23109 5859 23167 5865
rect 6273 5831 6331 5837
rect 6273 5797 6285 5831
rect 6319 5797 6331 5831
rect 6656 5828 6684 5856
rect 8018 5828 8024 5840
rect 6656 5800 8024 5828
rect 6273 5791 6331 5797
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 7064 5732 7113 5760
rect 7064 5720 7070 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7558 5760 7564 5772
rect 7519 5732 7564 5760
rect 7101 5723 7159 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7668 5769 7696 5800
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 13446 5788 13452 5840
rect 13504 5788 13510 5840
rect 16942 5788 16948 5840
rect 17000 5828 17006 5840
rect 17037 5831 17095 5837
rect 17037 5828 17049 5831
rect 17000 5800 17049 5828
rect 17000 5788 17006 5800
rect 17037 5797 17049 5800
rect 17083 5828 17095 5831
rect 17405 5831 17463 5837
rect 17405 5828 17417 5831
rect 17083 5800 17417 5828
rect 17083 5797 17095 5800
rect 17037 5791 17095 5797
rect 17405 5797 17417 5800
rect 17451 5828 17463 5831
rect 18230 5828 18236 5840
rect 17451 5800 18236 5828
rect 17451 5797 17463 5800
rect 17405 5791 17463 5797
rect 18230 5788 18236 5800
rect 18288 5788 18294 5840
rect 19886 5828 19892 5840
rect 19847 5800 19892 5828
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 22002 5788 22008 5840
rect 22060 5828 22066 5840
rect 22060 5800 22692 5828
rect 22060 5788 22066 5800
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5729 7711 5763
rect 9950 5760 9956 5772
rect 9911 5732 9956 5760
rect 7653 5723 7711 5729
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10468 5732 11345 5760
rect 10468 5720 10474 5732
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 11698 5760 11704 5772
rect 11379 5732 11704 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 12986 5760 12992 5772
rect 12947 5732 12992 5760
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13136 5732 13737 5760
rect 13136 5720 13142 5732
rect 13725 5729 13737 5732
rect 13771 5760 13783 5763
rect 14090 5760 14096 5772
rect 13771 5732 14096 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 19058 5760 19064 5772
rect 19019 5732 19064 5760
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 21818 5760 21824 5772
rect 20496 5732 21824 5760
rect 20496 5720 20502 5732
rect 21818 5720 21824 5732
rect 21876 5760 21882 5772
rect 22664 5769 22692 5800
rect 22281 5763 22339 5769
rect 22281 5760 22293 5763
rect 21876 5732 22293 5760
rect 21876 5720 21882 5732
rect 22281 5729 22293 5732
rect 22327 5729 22339 5763
rect 22281 5723 22339 5729
rect 22649 5763 22707 5769
rect 22649 5729 22661 5763
rect 22695 5729 22707 5763
rect 22830 5760 22836 5772
rect 22791 5732 22836 5760
rect 22649 5723 22707 5729
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 3436 5664 4261 5692
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4614 5692 4620 5704
rect 4571 5664 4620 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4264 5556 4292 5655
rect 4614 5652 4620 5664
rect 4672 5692 4678 5704
rect 5810 5692 5816 5704
rect 4672 5664 5816 5692
rect 4672 5652 4678 5664
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 8021 5627 8079 5633
rect 8021 5624 8033 5627
rect 7800 5596 8033 5624
rect 7800 5584 7806 5596
rect 8021 5593 8033 5596
rect 8067 5593 8079 5627
rect 8021 5587 8079 5593
rect 11238 5584 11244 5636
rect 11296 5624 11302 5636
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 11296 5596 11529 5624
rect 11296 5584 11302 5596
rect 11517 5593 11529 5596
rect 11563 5624 11575 5627
rect 13538 5624 13544 5636
rect 11563 5596 13544 5624
rect 11563 5593 11575 5596
rect 11517 5587 11575 5593
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 18141 5627 18199 5633
rect 18141 5593 18153 5627
rect 18187 5624 18199 5627
rect 18966 5624 18972 5636
rect 18187 5596 18972 5624
rect 18187 5593 18199 5596
rect 18141 5587 18199 5593
rect 18966 5584 18972 5596
rect 19024 5584 19030 5636
rect 21450 5584 21456 5636
rect 21508 5624 21514 5636
rect 22388 5624 22416 5655
rect 23566 5624 23572 5636
rect 21508 5596 23572 5624
rect 21508 5584 21514 5596
rect 23566 5584 23572 5596
rect 23624 5584 23630 5636
rect 4706 5556 4712 5568
rect 4264 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 8570 5556 8576 5568
rect 7156 5528 8576 5556
rect 7156 5516 7162 5528
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14148 5528 14749 5556
rect 14148 5516 14154 5528
rect 14737 5525 14749 5528
rect 14783 5556 14795 5559
rect 15470 5556 15476 5568
rect 14783 5528 15476 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 21361 5559 21419 5565
rect 21361 5525 21373 5559
rect 21407 5556 21419 5559
rect 22830 5556 22836 5568
rect 21407 5528 22836 5556
rect 21407 5525 21419 5528
rect 21361 5519 21419 5525
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 1104 5466 24656 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 24656 5466
rect 1104 5392 24656 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4982 5352 4988 5364
rect 4571 5324 4988 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5350 5352 5356 5364
rect 5311 5324 5356 5352
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 7558 5352 7564 5364
rect 6503 5324 7564 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 13078 5352 13084 5364
rect 12759 5324 13084 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 21450 5352 21456 5364
rect 21411 5324 21456 5352
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 22002 5352 22008 5364
rect 21963 5324 22008 5352
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 4157 5287 4215 5293
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4614 5284 4620 5296
rect 4203 5256 4620 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 4764 5256 4813 5284
rect 4764 5244 4770 5256
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 4801 5247 4859 5253
rect 6089 5287 6147 5293
rect 6089 5253 6101 5287
rect 6135 5284 6147 5287
rect 6638 5284 6644 5296
rect 6135 5256 6644 5284
rect 6135 5253 6147 5256
rect 6089 5247 6147 5253
rect 1670 5148 1676 5160
rect 1631 5120 1676 5148
rect 1670 5108 1676 5120
rect 1728 5108 1734 5160
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 2096 5120 2237 5148
rect 2096 5108 2102 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 4816 5148 4844 5247
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 12986 5244 12992 5296
rect 13044 5284 13050 5296
rect 13909 5287 13967 5293
rect 13909 5284 13921 5287
rect 13044 5256 13921 5284
rect 13044 5244 13050 5256
rect 13909 5253 13921 5256
rect 13955 5253 13967 5287
rect 13909 5247 13967 5253
rect 21085 5287 21143 5293
rect 21085 5253 21097 5287
rect 21131 5284 21143 5287
rect 22020 5284 22048 5312
rect 21131 5256 22048 5284
rect 21131 5253 21143 5256
rect 21085 5247 21143 5253
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6914 5216 6920 5228
rect 5767 5188 6920 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7742 5216 7748 5228
rect 7239 5188 7748 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 8812 5188 9505 5216
rect 8812 5176 8818 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 17681 5219 17739 5225
rect 15528 5188 16712 5216
rect 15528 5176 15534 5188
rect 7466 5148 7472 5160
rect 4816 5120 7472 5148
rect 2225 5111 2283 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8846 5108 8852 5160
rect 8904 5108 8910 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 10919 5120 11376 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 2590 5040 2596 5092
rect 2648 5040 2654 5092
rect 11348 5024 11376 5120
rect 11698 5108 11704 5160
rect 11756 5148 11762 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 11756 5120 13093 5148
rect 11756 5108 11762 5120
rect 13081 5117 13093 5120
rect 13127 5148 13139 5151
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 13127 5120 13553 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 13541 5117 13553 5120
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 16684 5157 16712 5188
rect 17681 5185 17693 5219
rect 17727 5216 17739 5219
rect 18509 5219 18567 5225
rect 18509 5216 18521 5219
rect 17727 5188 18521 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 18509 5185 18521 5188
rect 18555 5216 18567 5219
rect 19242 5216 19248 5228
rect 18555 5188 19248 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 19576 5188 20269 5216
rect 19576 5176 19582 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 15105 5151 15163 5157
rect 15105 5148 15117 5151
rect 14608 5120 15117 5148
rect 14608 5108 14614 5120
rect 15105 5117 15117 5120
rect 15151 5148 15163 5151
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 15151 5120 16221 5148
rect 15151 5117 15163 5120
rect 15105 5111 15163 5117
rect 16209 5117 16221 5120
rect 16255 5117 16267 5151
rect 16209 5111 16267 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 16715 5120 17141 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 17129 5117 17141 5120
rect 17175 5148 17187 5151
rect 17586 5148 17592 5160
rect 17175 5120 17592 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 18230 5148 18236 5160
rect 18191 5120 18236 5148
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 21818 5148 21824 5160
rect 21779 5120 21824 5148
rect 21818 5108 21824 5120
rect 21876 5148 21882 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 21876 5120 22753 5148
rect 21876 5108 21882 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 14090 5080 14096 5092
rect 13372 5052 14096 5080
rect 9950 4972 9956 5024
rect 10008 5012 10014 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 10008 4984 10057 5012
rect 10008 4972 10014 4984
rect 10045 4981 10057 4984
rect 10091 5012 10103 5015
rect 10870 5012 10876 5024
rect 10091 4984 10876 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 13265 5015 13323 5021
rect 13265 4981 13277 5015
rect 13311 5012 13323 5015
rect 13372 5012 13400 5052
rect 14090 5040 14096 5052
rect 14148 5040 14154 5092
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 14461 5083 14519 5089
rect 14461 5080 14473 5083
rect 14240 5052 14473 5080
rect 14240 5040 14246 5052
rect 14461 5049 14473 5052
rect 14507 5049 14519 5083
rect 14461 5043 14519 5049
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 16114 5080 16120 5092
rect 15611 5052 16120 5080
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 16114 5040 16120 5052
rect 16172 5040 16178 5092
rect 18966 5040 18972 5092
rect 19024 5040 19030 5092
rect 15838 5012 15844 5024
rect 13311 4984 13400 5012
rect 15799 4984 15844 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 16850 5012 16856 5024
rect 16811 4984 16856 5012
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 1104 4922 24656 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 24656 4922
rect 1104 4848 24656 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4808 2102 4820
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 2096 4780 2329 4808
rect 2096 4768 2102 4780
rect 2317 4777 2329 4780
rect 2363 4777 2375 4811
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 2317 4771 2375 4777
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 3602 4808 3608 4820
rect 3467 4780 3608 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 4890 4808 4896 4820
rect 4847 4780 4896 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4816 4672 4844 4771
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 8846 4808 8852 4820
rect 7883 4780 8852 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12216 4780 12357 4808
rect 12216 4768 12222 4780
rect 12345 4777 12357 4780
rect 12391 4808 12403 4811
rect 13630 4808 13636 4820
rect 12391 4780 13636 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 13630 4768 13636 4780
rect 13688 4808 13694 4820
rect 18417 4811 18475 4817
rect 13688 4780 13814 4808
rect 13688 4768 13694 4780
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 5776 4712 6408 4740
rect 5776 4700 5782 4712
rect 4295 4644 4844 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 5408 4644 5917 4672
rect 5408 4632 5414 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6380 4681 6408 4712
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 8110 4740 8116 4752
rect 7524 4712 8116 4740
rect 7524 4700 7530 4712
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 13538 4740 13544 4752
rect 13499 4712 13544 4740
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 6365 4675 6423 4681
rect 6052 4644 6097 4672
rect 6052 4632 6058 4644
rect 6365 4641 6377 4675
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 8570 4672 8576 4684
rect 6512 4644 6557 4672
rect 8531 4644 8576 4672
rect 6512 4632 6518 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 9858 4672 9864 4684
rect 9771 4644 9864 4672
rect 9858 4632 9864 4644
rect 9916 4672 9922 4684
rect 11146 4672 11152 4684
rect 9916 4644 11152 4672
rect 9916 4632 9922 4644
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 12989 4675 13047 4681
rect 12989 4641 13001 4675
rect 13035 4672 13047 4675
rect 13556 4672 13584 4700
rect 13035 4644 13584 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 7055 4576 7389 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7377 4573 7389 4576
rect 7423 4604 7435 4607
rect 7466 4604 7472 4616
rect 7423 4576 7472 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 13786 4604 13814 4780
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 18966 4808 18972 4820
rect 18463 4780 18972 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 20864 4780 21373 4808
rect 20864 4768 20870 4780
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 21361 4771 21419 4777
rect 21818 4768 21824 4820
rect 21876 4808 21882 4820
rect 22005 4811 22063 4817
rect 22005 4808 22017 4811
rect 21876 4780 22017 4808
rect 21876 4768 21882 4780
rect 22005 4777 22017 4780
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 18785 4743 18843 4749
rect 18785 4709 18797 4743
rect 18831 4740 18843 4743
rect 19610 4740 19616 4752
rect 18831 4712 19616 4740
rect 18831 4709 18843 4712
rect 18785 4703 18843 4709
rect 19610 4700 19616 4712
rect 19668 4740 19674 4752
rect 19978 4740 19984 4752
rect 19668 4712 19984 4740
rect 19668 4700 19674 4712
rect 19978 4700 19984 4712
rect 20036 4700 20042 4752
rect 21729 4743 21787 4749
rect 21729 4709 21741 4743
rect 21775 4740 21787 4743
rect 22830 4740 22836 4752
rect 21775 4712 22836 4740
rect 21775 4709 21787 4712
rect 21729 4703 21787 4709
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 16850 4632 16856 4684
rect 16908 4632 16914 4684
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 17644 4644 18245 4672
rect 17644 4632 17650 4644
rect 18233 4641 18245 4644
rect 18279 4672 18291 4675
rect 19058 4672 19064 4684
rect 18279 4644 19064 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 21177 4675 21235 4681
rect 21177 4672 21189 4675
rect 19484 4644 21189 4672
rect 19484 4632 19490 4644
rect 21177 4641 21189 4644
rect 21223 4672 21235 4675
rect 22462 4672 22468 4684
rect 21223 4644 22468 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4672 23535 4675
rect 23566 4672 23572 4684
rect 23523 4644 23572 4672
rect 23523 4641 23535 4644
rect 23477 4635 23535 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 13786 4576 14565 4604
rect 14553 4573 14565 4576
rect 14599 4604 14611 4607
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 14599 4576 15485 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15746 4604 15752 4616
rect 15707 4576 15752 4604
rect 15473 4567 15531 4573
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 10045 4539 10103 4545
rect 10045 4536 10057 4539
rect 8536 4508 10057 4536
rect 8536 4496 8542 4508
rect 10045 4505 10057 4508
rect 10091 4505 10103 4539
rect 10045 4499 10103 4505
rect 11517 4539 11575 4545
rect 11517 4505 11529 4539
rect 11563 4536 11575 4539
rect 12618 4536 12624 4548
rect 11563 4508 12624 4536
rect 11563 4505 11575 4508
rect 11517 4499 11575 4505
rect 12618 4496 12624 4508
rect 12676 4496 12682 4548
rect 14274 4496 14280 4548
rect 14332 4536 14338 4548
rect 14829 4539 14887 4545
rect 14829 4536 14841 4539
rect 14332 4508 14841 4536
rect 14332 4496 14338 4508
rect 14829 4505 14841 4508
rect 14875 4505 14887 4539
rect 14829 4499 14887 4505
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 4433 4471 4491 4477
rect 4433 4468 4445 4471
rect 3752 4440 4445 4468
rect 3752 4428 3758 4440
rect 4433 4437 4445 4440
rect 4479 4437 4491 4471
rect 5350 4468 5356 4480
rect 5311 4440 5356 4468
rect 4433 4431 4491 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 6972 4440 8769 4468
rect 6972 4428 6978 4440
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 12713 4471 12771 4477
rect 12713 4437 12725 4471
rect 12759 4468 12771 4471
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 12759 4440 13185 4468
rect 12759 4437 12771 4440
rect 12713 4431 12771 4437
rect 13173 4437 13185 4440
rect 13219 4468 13231 4471
rect 13354 4468 13360 4480
rect 13219 4440 13360 4468
rect 13219 4437 13231 4440
rect 13173 4431 13231 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 15488 4468 15516 4567
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 16298 4564 16304 4616
rect 16356 4604 16362 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16356 4576 17509 4604
rect 16356 4564 16362 4576
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 21634 4564 21640 4616
rect 21692 4604 21698 4616
rect 22373 4607 22431 4613
rect 22373 4604 22385 4607
rect 21692 4576 22385 4604
rect 21692 4564 21698 4576
rect 22373 4573 22385 4576
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 16942 4468 16948 4480
rect 15488 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17954 4468 17960 4480
rect 17915 4440 17960 4468
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 20165 4471 20223 4477
rect 20165 4468 20177 4471
rect 20036 4440 20177 4468
rect 20036 4428 20042 4440
rect 20165 4437 20177 4440
rect 20211 4437 20223 4471
rect 20165 4431 20223 4437
rect 20533 4471 20591 4477
rect 20533 4437 20545 4471
rect 20579 4468 20591 4471
rect 20622 4468 20628 4480
rect 20579 4440 20628 4468
rect 20579 4437 20591 4440
rect 20533 4431 20591 4437
rect 20622 4428 20628 4440
rect 20680 4468 20686 4480
rect 21910 4468 21916 4480
rect 20680 4440 21916 4468
rect 20680 4428 20686 4440
rect 21910 4428 21916 4440
rect 21968 4428 21974 4480
rect 1104 4378 24656 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 24656 4378
rect 1104 4304 24656 4326
rect 2590 4264 2596 4276
rect 2551 4236 2596 4264
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5534 4264 5540 4276
rect 5491 4236 5540 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 6454 4264 6460 4276
rect 5592 4236 6460 4264
rect 5592 4224 5598 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7282 4264 7288 4276
rect 7208 4236 7288 4264
rect 2608 4196 2636 4224
rect 2608 4168 2728 4196
rect 2700 4128 2728 4168
rect 4798 4156 4804 4208
rect 4856 4196 4862 4208
rect 5350 4196 5356 4208
rect 4856 4168 5356 4196
rect 4856 4156 4862 4168
rect 5350 4156 5356 4168
rect 5408 4196 5414 4208
rect 7098 4196 7104 4208
rect 5408 4168 7104 4196
rect 5408 4156 5414 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 7208 4137 7236 4236
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 9769 4267 9827 4273
rect 9769 4233 9781 4267
rect 9815 4264 9827 4267
rect 9858 4264 9864 4276
rect 9815 4236 9864 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 10870 4264 10876 4276
rect 10831 4236 10876 4264
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17129 4267 17187 4273
rect 17129 4264 17141 4267
rect 16908 4236 17141 4264
rect 16908 4224 16914 4236
rect 17129 4233 17141 4236
rect 17175 4233 17187 4267
rect 17586 4264 17592 4276
rect 17547 4236 17592 4264
rect 17129 4227 17187 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 22462 4264 22468 4276
rect 22423 4236 22468 4264
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 22925 4267 22983 4273
rect 22925 4233 22937 4267
rect 22971 4264 22983 4267
rect 23566 4264 23572 4276
rect 22971 4236 23572 4264
rect 22971 4233 22983 4236
rect 22925 4227 22983 4233
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 15197 4199 15255 4205
rect 15197 4165 15209 4199
rect 15243 4196 15255 4199
rect 15746 4196 15752 4208
rect 15243 4168 15752 4196
rect 15243 4165 15255 4168
rect 15197 4159 15255 4165
rect 15746 4156 15752 4168
rect 15804 4196 15810 4208
rect 16577 4199 16635 4205
rect 16577 4196 16589 4199
rect 15804 4168 16589 4196
rect 15804 4156 15810 4168
rect 16577 4165 16589 4168
rect 16623 4165 16635 4199
rect 16577 4159 16635 4165
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2700 4100 3249 4128
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7193 4091 7251 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12216 4100 12633 4128
rect 12216 4088 12222 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12894 4128 12900 4140
rect 12807 4100 12900 4128
rect 12621 4091 12679 4097
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 13446 4128 13452 4140
rect 12952 4100 13452 4128
rect 12952 4088 12958 4100
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14550 4128 14556 4140
rect 13964 4100 14556 4128
rect 13964 4088 13970 4100
rect 14550 4088 14556 4100
rect 14608 4128 14614 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14608 4100 14657 4128
rect 14608 4088 14614 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 14792 4100 15700 4128
rect 14792 4088 14798 4100
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4029 3019 4063
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 2961 4023 3019 4029
rect 10244 4032 10609 4060
rect 2976 3992 3004 4023
rect 3142 3992 3148 4004
rect 2976 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3694 3952 3700 4004
rect 3752 3952 3758 4004
rect 4985 3995 5043 4001
rect 4985 3961 4997 3995
rect 5031 3992 5043 3995
rect 5442 3992 5448 4004
rect 5031 3964 5448 3992
rect 5031 3961 5043 3964
rect 4985 3955 5043 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6457 3995 6515 4001
rect 6457 3961 6469 3995
rect 6503 3992 6515 3995
rect 9214 3992 9220 4004
rect 6503 3964 7972 3992
rect 9175 3964 9220 3992
rect 6503 3961 6515 3964
rect 6457 3955 6515 3961
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7944 3924 7972 3964
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 8478 3924 8484 3936
rect 7944 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 10244 3933 10272 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 10735 4032 11560 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 11532 4001 11560 4032
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 15470 4060 15476 4072
rect 14332 4032 15476 4060
rect 14332 4020 14338 4032
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15672 4069 15700 4100
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 21910 4128 21916 4140
rect 20036 4100 21772 4128
rect 21871 4100 21916 4128
rect 20036 4088 20042 4100
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 15838 4060 15844 4072
rect 15703 4032 15844 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 16114 4060 16120 4072
rect 16075 4032 16120 4060
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 11517 3995 11575 4001
rect 11517 3961 11529 3995
rect 11563 3992 11575 3995
rect 11563 3964 12020 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9640 3896 10241 3924
rect 9640 3884 9646 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11388 3896 11805 3924
rect 11388 3884 11394 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11992 3924 12020 3964
rect 13354 3952 13360 4004
rect 13412 3952 13418 4004
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 14918 3992 14924 4004
rect 14240 3964 14924 3992
rect 14240 3952 14246 3964
rect 14918 3952 14924 3964
rect 14976 3992 14982 4004
rect 16224 3992 16252 4023
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18012 4032 19165 4060
rect 18012 4020 18018 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19610 4060 19616 4072
rect 19523 4032 19616 4060
rect 19153 4023 19211 4029
rect 14976 3964 16252 3992
rect 14976 3952 14982 3964
rect 17402 3924 17408 3936
rect 11992 3896 17408 3924
rect 11793 3887 11851 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 19168 3924 19196 4023
rect 19610 4020 19616 4032
rect 19668 4060 19674 4072
rect 20346 4060 20352 4072
rect 19668 4032 20352 4060
rect 19668 4020 19674 4032
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 21450 4060 21456 4072
rect 20763 4032 21456 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 21634 4060 21640 4072
rect 21547 4032 21640 4060
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 21744 4060 21772 4100
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 22002 4060 22008 4072
rect 21744 4032 22008 4060
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 19242 3952 19248 4004
rect 19300 3952 19306 4004
rect 20898 3952 20904 4004
rect 20956 3992 20962 4004
rect 21652 3992 21680 4020
rect 20956 3964 21680 3992
rect 20956 3952 20962 3964
rect 20438 3924 20444 3936
rect 19168 3896 20444 3924
rect 20438 3884 20444 3896
rect 20496 3924 20502 3936
rect 21269 3927 21327 3933
rect 21269 3924 21281 3927
rect 20496 3896 21281 3924
rect 20496 3884 20502 3896
rect 21269 3893 21281 3896
rect 21315 3924 21327 3927
rect 22646 3924 22652 3936
rect 21315 3896 22652 3924
rect 21315 3893 21327 3896
rect 21269 3887 21327 3893
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 1104 3834 24656 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 24656 3834
rect 1104 3760 24656 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3694 3720 3700 3732
rect 3099 3692 3700 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 4798 3720 4804 3732
rect 4759 3692 4804 3720
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 12713 3723 12771 3729
rect 12713 3689 12725 3723
rect 12759 3720 12771 3723
rect 12894 3720 12900 3732
rect 12759 3692 12900 3720
rect 12759 3689 12771 3692
rect 12713 3683 12771 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14918 3720 14924 3732
rect 14879 3692 14924 3720
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 20027 3692 21864 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 21836 3664 21864 3692
rect 5442 3652 5448 3664
rect 5184 3624 5448 3652
rect 5184 3593 5212 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 8527 3624 10517 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 10505 3621 10517 3624
rect 10551 3652 10563 3655
rect 10594 3652 10600 3664
rect 10551 3624 10600 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 11514 3612 11520 3664
rect 11572 3612 11578 3664
rect 12253 3655 12311 3661
rect 12253 3621 12265 3655
rect 12299 3652 12311 3655
rect 14550 3652 14556 3664
rect 12299 3624 14556 3652
rect 12299 3621 12311 3624
rect 12253 3615 12311 3621
rect 14550 3612 14556 3624
rect 14608 3612 14614 3664
rect 16114 3652 16120 3664
rect 15212 3624 16120 3652
rect 3697 3587 3755 3593
rect 3697 3553 3709 3587
rect 3743 3584 3755 3587
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 3743 3556 5181 3584
rect 3743 3553 3755 3556
rect 3697 3547 3755 3553
rect 5169 3553 5181 3556
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 5534 3584 5540 3596
rect 5316 3556 5540 3584
rect 5316 3544 5322 3556
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6052 3556 6653 3584
rect 6052 3544 6058 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 7156 3556 7205 3584
rect 7156 3544 7162 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 13817 3587 13875 3593
rect 13817 3584 13829 3587
rect 11940 3556 13829 3584
rect 11940 3544 11946 3556
rect 13817 3553 13829 3556
rect 13863 3584 13875 3587
rect 13906 3584 13912 3596
rect 13863 3556 13912 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14182 3584 14188 3596
rect 14143 3556 14188 3584
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 15212 3584 15240 3624
rect 16114 3612 16120 3624
rect 16172 3652 16178 3664
rect 16209 3655 16267 3661
rect 16209 3652 16221 3655
rect 16172 3624 16221 3652
rect 16172 3612 16178 3624
rect 16209 3621 16221 3624
rect 16255 3621 16267 3655
rect 16209 3615 16267 3621
rect 17678 3612 17684 3664
rect 17736 3612 17742 3664
rect 21818 3612 21824 3664
rect 21876 3612 21882 3664
rect 14415 3556 15240 3584
rect 16025 3587 16083 3593
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 16025 3553 16037 3587
rect 16071 3584 16083 3587
rect 16298 3584 16304 3596
rect 16071 3556 16304 3584
rect 16071 3553 16083 3556
rect 16025 3547 16083 3553
rect 4982 3516 4988 3528
rect 4943 3488 4988 3516
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14384 3516 14412 3547
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 16942 3584 16948 3596
rect 16903 3556 16948 3584
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 19797 3587 19855 3593
rect 19797 3584 19809 3587
rect 19116 3556 19809 3584
rect 19116 3544 19122 3556
rect 19797 3553 19809 3556
rect 19843 3584 19855 3587
rect 20257 3587 20315 3593
rect 20257 3584 20269 3587
rect 19843 3556 20269 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 20257 3553 20269 3556
rect 20303 3553 20315 3587
rect 20257 3547 20315 3553
rect 17218 3516 17224 3528
rect 13780 3488 14412 3516
rect 17179 3488 17224 3516
rect 13780 3476 13786 3488
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 18966 3516 18972 3528
rect 18927 3488 18972 3516
rect 18966 3476 18972 3488
rect 19024 3516 19030 3528
rect 20898 3516 20904 3528
rect 19024 3488 20904 3516
rect 19024 3476 19030 3488
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 21082 3516 21088 3528
rect 21043 3488 21088 3516
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 23109 3519 23167 3525
rect 23109 3516 23121 3519
rect 21508 3488 23121 3516
rect 21508 3476 21514 3488
rect 23109 3485 23121 3488
rect 23155 3485 23167 3519
rect 23109 3479 23167 3485
rect 5994 3380 6000 3392
rect 5955 3352 6000 3380
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 8846 3380 8852 3392
rect 8628 3352 8852 3380
rect 8628 3340 8634 3352
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 13449 3383 13507 3389
rect 13449 3349 13461 3383
rect 13495 3380 13507 3383
rect 14734 3380 14740 3392
rect 13495 3352 14740 3380
rect 13495 3349 13507 3352
rect 13449 3343 13507 3349
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 19521 3383 19579 3389
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 19978 3380 19984 3392
rect 19567 3352 19984 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 1104 3290 24656 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 24656 3290
rect 1104 3216 24656 3238
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 8904 3148 9873 3176
rect 8904 3136 8910 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 10919 3148 11437 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 11425 3145 11437 3148
rect 11471 3176 11483 3179
rect 11514 3176 11520 3188
rect 11471 3148 11520 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12894 3176 12900 3188
rect 12855 3148 12900 3176
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13541 3179 13599 3185
rect 13541 3145 13553 3179
rect 13587 3176 13599 3179
rect 13630 3176 13636 3188
rect 13587 3148 13636 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 13630 3136 13636 3148
rect 13688 3176 13694 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 13688 3148 16129 3176
rect 13688 3136 13694 3148
rect 16117 3145 16129 3148
rect 16163 3176 16175 3179
rect 16298 3176 16304 3188
rect 16163 3148 16304 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16669 3179 16727 3185
rect 16669 3145 16681 3179
rect 16715 3176 16727 3179
rect 16942 3176 16948 3188
rect 16715 3148 16948 3176
rect 16715 3145 16727 3148
rect 16669 3139 16727 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 17678 3176 17684 3188
rect 17451 3148 17684 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 20346 3176 20352 3188
rect 20259 3148 20352 3176
rect 20346 3136 20352 3148
rect 20404 3176 20410 3188
rect 20404 3148 21680 3176
rect 20404 3136 20410 3148
rect 8110 3108 8116 3120
rect 2056 3080 7972 3108
rect 8023 3080 8116 3108
rect 2056 3052 2084 3080
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 2038 3040 2044 3052
rect 1636 3012 2044 3040
rect 1636 3000 1642 3012
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 5718 3040 5724 3052
rect 4663 3012 5724 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 5718 3000 5724 3012
rect 5776 3040 5782 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 5776 3012 7021 3040
rect 5776 3000 5782 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7944 3040 7972 3080
rect 8110 3068 8116 3080
rect 8168 3108 8174 3120
rect 10226 3108 10232 3120
rect 8168 3080 10232 3108
rect 8168 3068 8174 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 7944 3012 9321 3040
rect 7009 3003 7067 3009
rect 9309 3009 9321 3012
rect 9355 3040 9367 3043
rect 9582 3040 9588 3052
rect 9355 3012 9588 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 15749 3043 15807 3049
rect 11992 3012 12756 3040
rect 11992 2984 12020 3012
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2941 2191 2975
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 2133 2935 2191 2941
rect 3068 2944 3525 2972
rect 2148 2904 2176 2935
rect 2590 2904 2596 2916
rect 1688 2876 2176 2904
rect 2551 2876 2596 2904
rect 290 2796 296 2848
rect 348 2836 354 2848
rect 1688 2845 1716 2876
rect 2590 2864 2596 2876
rect 2648 2864 2654 2916
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 348 2808 1685 2836
rect 348 2796 354 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 3068 2845 3096 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 5442 2972 5448 2984
rect 4203 2944 5304 2972
rect 5403 2944 5448 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 5166 2904 5172 2916
rect 5127 2876 5172 2904
rect 5166 2864 5172 2876
rect 5224 2864 5230 2916
rect 5276 2904 5304 2944
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 7653 2975 7711 2981
rect 7653 2972 7665 2975
rect 7616 2944 7665 2972
rect 7616 2932 7622 2944
rect 7653 2941 7665 2944
rect 7699 2972 7711 2975
rect 9214 2972 9220 2984
rect 7699 2944 9220 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 11238 2972 11244 2984
rect 9723 2944 10548 2972
rect 11199 2944 11244 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 9766 2904 9772 2916
rect 5276 2876 9772 2904
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 10520 2913 10548 2944
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11974 2972 11980 2984
rect 11935 2944 11980 2972
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 12618 2972 12624 2984
rect 12579 2944 12624 2972
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 12728 2981 12756 3012
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 15795 3012 16957 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 16945 3009 16957 3012
rect 16991 3040 17003 3043
rect 17218 3040 17224 3052
rect 16991 3012 17224 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 19426 3040 19432 3052
rect 19387 3012 19432 3040
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 20364 3049 20392 3136
rect 21358 3108 21364 3120
rect 21319 3080 21364 3108
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 21652 3108 21680 3148
rect 21818 3136 21824 3188
rect 21876 3176 21882 3188
rect 21913 3179 21971 3185
rect 21913 3176 21925 3179
rect 21876 3148 21925 3176
rect 21876 3136 21882 3148
rect 21913 3145 21925 3148
rect 21959 3145 21971 3179
rect 22646 3176 22652 3188
rect 22607 3148 22652 3176
rect 21913 3139 21971 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 22281 3111 22339 3117
rect 22281 3108 22293 3111
rect 21652 3080 22293 3108
rect 22281 3077 22293 3080
rect 22327 3077 22339 3111
rect 22281 3071 22339 3077
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 12713 2935 12771 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15470 2972 15476 2984
rect 15243 2944 15476 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 18524 2944 18889 2972
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 12066 2904 12072 2916
rect 10551 2876 12072 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2740 2808 3065 2836
rect 2740 2796 2746 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5994 2836 6000 2848
rect 4764 2808 6000 2836
rect 4764 2796 4770 2808
rect 5994 2796 6000 2808
rect 6052 2836 6058 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6052 2808 6377 2836
rect 6052 2796 6058 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 11330 2836 11336 2848
rect 10192 2808 11336 2836
rect 10192 2796 10198 2808
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 15286 2836 15292 2848
rect 14424 2808 15292 2836
rect 14424 2796 14430 2808
rect 15286 2796 15292 2808
rect 15344 2836 15350 2848
rect 18524 2845 18552 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 18969 2975 19027 2981
rect 18969 2941 18981 2975
rect 19015 2972 19027 2975
rect 20438 2972 20444 2984
rect 19015 2944 19840 2972
rect 20399 2944 20444 2972
rect 19015 2941 19027 2944
rect 18969 2935 19027 2941
rect 19812 2913 19840 2944
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 20907 2975 20965 2981
rect 20907 2972 20919 2975
rect 20680 2944 20919 2972
rect 20680 2932 20686 2944
rect 20907 2941 20919 2944
rect 20953 2941 20965 2975
rect 20907 2935 20965 2941
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2972 21051 2975
rect 22002 2972 22008 2984
rect 21039 2944 22008 2972
rect 21039 2941 21051 2944
rect 20993 2935 21051 2941
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 19797 2907 19855 2913
rect 19797 2873 19809 2907
rect 19843 2904 19855 2907
rect 19886 2904 19892 2916
rect 19843 2876 19892 2904
rect 19843 2873 19855 2876
rect 19797 2867 19855 2873
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 21082 2864 21088 2916
rect 21140 2904 21146 2916
rect 23017 2907 23075 2913
rect 23017 2904 23029 2907
rect 21140 2876 23029 2904
rect 21140 2864 21146 2876
rect 23017 2873 23029 2876
rect 23063 2873 23075 2907
rect 23017 2867 23075 2873
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 15344 2808 18521 2836
rect 15344 2796 15350 2808
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 1104 2746 24656 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 24656 2746
rect 1104 2672 24656 2694
rect 2038 2632 2044 2644
rect 1999 2604 2044 2632
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 3605 2635 3663 2641
rect 3605 2632 3617 2635
rect 2648 2604 3617 2632
rect 2648 2592 2654 2604
rect 3605 2601 3617 2604
rect 3651 2632 3663 2635
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 3651 2604 4169 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4706 2632 4712 2644
rect 4479 2604 4712 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5166 2632 5172 2644
rect 4847 2604 5172 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10594 2632 10600 2644
rect 10555 2604 10600 2632
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11238 2632 11244 2644
rect 11199 2604 11244 2632
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12676 2604 13277 2632
rect 12676 2592 12682 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13722 2632 13728 2644
rect 13683 2604 13728 2632
rect 13265 2595 13323 2601
rect 4982 2524 4988 2576
rect 5040 2564 5046 2576
rect 5077 2567 5135 2573
rect 5077 2564 5089 2567
rect 5040 2536 5089 2564
rect 5040 2524 5046 2536
rect 5077 2533 5089 2536
rect 5123 2564 5135 2567
rect 7576 2564 7604 2592
rect 5123 2536 7604 2564
rect 13280 2564 13308 2595
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14182 2632 14188 2644
rect 14139 2604 14188 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 15470 2632 15476 2644
rect 14507 2604 15476 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 14366 2564 14372 2576
rect 13280 2536 14372 2564
rect 5123 2533 5135 2536
rect 5077 2527 5135 2533
rect 14366 2524 14372 2536
rect 14424 2524 14430 2576
rect 12253 2499 12311 2505
rect 12253 2465 12265 2499
rect 12299 2496 12311 2499
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 12299 2468 12817 2496
rect 12299 2465 12311 2468
rect 12253 2459 12311 2465
rect 12805 2465 12817 2468
rect 12851 2496 12863 2499
rect 12894 2496 12900 2508
rect 12851 2468 12900 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 12989 2363 13047 2369
rect 12989 2329 13001 2363
rect 13035 2360 13047 2363
rect 14476 2360 14504 2595
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 17736 2604 18705 2632
rect 17736 2592 17742 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 19058 2632 19064 2644
rect 19019 2604 19064 2632
rect 18693 2595 18751 2601
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19978 2632 19984 2644
rect 19939 2604 19984 2632
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20622 2632 20628 2644
rect 20583 2604 20628 2632
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 21358 2632 21364 2644
rect 21319 2604 21364 2632
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 21450 2592 21456 2644
rect 21508 2632 21514 2644
rect 21729 2635 21787 2641
rect 21729 2632 21741 2635
rect 21508 2604 21741 2632
rect 21508 2592 21514 2604
rect 21729 2601 21741 2604
rect 21775 2632 21787 2635
rect 21775 2604 22232 2632
rect 21775 2601 21787 2604
rect 21729 2595 21787 2601
rect 14734 2564 14740 2576
rect 14695 2536 14740 2564
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 19076 2496 19104 2592
rect 20640 2564 20668 2592
rect 22097 2567 22155 2573
rect 22097 2564 22109 2567
rect 20640 2536 22109 2564
rect 22097 2533 22109 2536
rect 22143 2533 22155 2567
rect 22097 2527 22155 2533
rect 22204 2505 22232 2604
rect 18555 2468 19104 2496
rect 19613 2499 19671 2505
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 19613 2465 19625 2499
rect 19659 2465 19671 2499
rect 19613 2459 19671 2465
rect 22189 2499 22247 2505
rect 22189 2465 22201 2499
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2428 18015 2431
rect 18966 2428 18972 2440
rect 18003 2400 18972 2428
rect 18003 2397 18015 2400
rect 17957 2391 18015 2397
rect 18966 2388 18972 2400
rect 19024 2428 19030 2440
rect 19628 2428 19656 2459
rect 19024 2400 19656 2428
rect 19024 2388 19030 2400
rect 13035 2332 14504 2360
rect 13035 2329 13047 2332
rect 12989 2323 13047 2329
rect 1104 2202 24656 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 24656 2202
rect 1104 2128 24656 2150
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 22370 1340 22376 1352
rect 12216 1312 22376 1340
rect 12216 1300 12222 1312
rect 22370 1300 22376 1312
rect 22428 1300 22434 1352
rect 4890 8 4896 60
rect 4948 48 4954 60
rect 15194 48 15200 60
rect 4948 20 15200 48
rect 4948 8 4954 20
rect 15194 8 15200 20
rect 15252 8 15258 60
<< via1 >>
rect 8392 27208 8444 27260
rect 11704 27208 11756 27260
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 4988 25347 5040 25356
rect 4988 25313 4997 25347
rect 4997 25313 5031 25347
rect 5031 25313 5040 25347
rect 4988 25304 5040 25313
rect 5540 25304 5592 25356
rect 8392 25347 8444 25356
rect 8392 25313 8401 25347
rect 8401 25313 8435 25347
rect 8435 25313 8444 25347
rect 8392 25304 8444 25313
rect 12624 25304 12676 25356
rect 13176 25304 13228 25356
rect 16120 25304 16172 25356
rect 16764 25347 16816 25356
rect 16764 25313 16773 25347
rect 16773 25313 16807 25347
rect 16807 25313 16816 25347
rect 16764 25304 16816 25313
rect 22468 25304 22520 25356
rect 2044 25236 2096 25288
rect 7288 25236 7340 25288
rect 14188 25168 14240 25220
rect 5172 25143 5224 25152
rect 5172 25109 5181 25143
rect 5181 25109 5215 25143
rect 5215 25109 5224 25143
rect 5172 25100 5224 25109
rect 8576 25143 8628 25152
rect 8576 25109 8585 25143
rect 8585 25109 8619 25143
rect 8619 25109 8628 25143
rect 8576 25100 8628 25109
rect 9404 25100 9456 25152
rect 10416 25100 10468 25152
rect 10876 25143 10928 25152
rect 10876 25109 10885 25143
rect 10885 25109 10919 25143
rect 10919 25109 10928 25143
rect 10876 25100 10928 25109
rect 13544 25100 13596 25152
rect 14464 25143 14516 25152
rect 14464 25109 14473 25143
rect 14473 25109 14507 25143
rect 14507 25109 14516 25143
rect 14464 25100 14516 25109
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 22560 25143 22612 25152
rect 22560 25109 22569 25143
rect 22569 25109 22603 25143
rect 22603 25109 22612 25143
rect 22560 25100 22612 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 4988 24896 5040 24948
rect 7288 24939 7340 24948
rect 7288 24905 7297 24939
rect 7297 24905 7331 24939
rect 7331 24905 7340 24939
rect 7288 24896 7340 24905
rect 8300 24939 8352 24948
rect 8300 24905 8309 24939
rect 8309 24905 8343 24939
rect 8343 24905 8352 24939
rect 8300 24896 8352 24905
rect 16120 24939 16172 24948
rect 16120 24905 16129 24939
rect 16129 24905 16163 24939
rect 16163 24905 16172 24939
rect 16120 24896 16172 24905
rect 16764 24939 16816 24948
rect 16764 24905 16773 24939
rect 16773 24905 16807 24939
rect 16807 24905 16816 24939
rect 16764 24896 16816 24905
rect 22468 24939 22520 24948
rect 22468 24905 22477 24939
rect 22477 24905 22511 24939
rect 22511 24905 22520 24939
rect 22468 24896 22520 24905
rect 23112 24939 23164 24948
rect 23112 24905 23121 24939
rect 23121 24905 23155 24939
rect 23155 24905 23164 24939
rect 23112 24896 23164 24905
rect 25504 24828 25556 24880
rect 9404 24803 9456 24812
rect 5172 24692 5224 24744
rect 6368 24692 6420 24744
rect 7288 24692 7340 24744
rect 7564 24692 7616 24744
rect 8024 24735 8076 24744
rect 8024 24701 8033 24735
rect 8033 24701 8067 24735
rect 8067 24701 8076 24735
rect 8024 24692 8076 24701
rect 9404 24769 9413 24803
rect 9413 24769 9447 24803
rect 9447 24769 9456 24803
rect 9404 24760 9456 24769
rect 10416 24760 10468 24812
rect 11060 24760 11112 24812
rect 13176 24803 13228 24812
rect 10600 24692 10652 24744
rect 10876 24735 10928 24744
rect 10876 24701 10885 24735
rect 10885 24701 10919 24735
rect 10919 24701 10928 24735
rect 10876 24692 10928 24701
rect 13176 24769 13185 24803
rect 13185 24769 13219 24803
rect 13219 24769 13228 24803
rect 13176 24760 13228 24769
rect 14188 24735 14240 24744
rect 9864 24624 9916 24676
rect 11520 24667 11572 24676
rect 11520 24633 11529 24667
rect 11529 24633 11563 24667
rect 11563 24633 11572 24667
rect 11520 24624 11572 24633
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 14464 24692 14516 24744
rect 15936 24692 15988 24744
rect 18880 24735 18932 24744
rect 18880 24701 18889 24735
rect 18889 24701 18923 24735
rect 18923 24701 18932 24735
rect 18880 24692 18932 24701
rect 18972 24692 19024 24744
rect 14924 24624 14976 24676
rect 4712 24556 4764 24608
rect 5356 24556 5408 24608
rect 8392 24556 8444 24608
rect 13084 24556 13136 24608
rect 17316 24599 17368 24608
rect 17316 24565 17325 24599
rect 17325 24565 17359 24599
rect 17359 24565 17368 24599
rect 17316 24556 17368 24565
rect 18696 24556 18748 24608
rect 21456 24692 21508 24744
rect 21732 24556 21784 24608
rect 23112 24692 23164 24744
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 8024 24352 8076 24404
rect 14188 24352 14240 24404
rect 15476 24352 15528 24404
rect 17316 24352 17368 24404
rect 3332 24284 3384 24336
rect 1676 24259 1728 24268
rect 1676 24225 1685 24259
rect 1685 24225 1719 24259
rect 1719 24225 1728 24259
rect 1676 24216 1728 24225
rect 4620 24259 4672 24268
rect 4620 24225 4629 24259
rect 4629 24225 4663 24259
rect 4663 24225 4672 24259
rect 4620 24216 4672 24225
rect 4712 24259 4764 24268
rect 4712 24225 4721 24259
rect 4721 24225 4755 24259
rect 4755 24225 4764 24259
rect 5172 24259 5224 24268
rect 4712 24216 4764 24225
rect 5172 24225 5181 24259
rect 5181 24225 5215 24259
rect 5215 24225 5224 24259
rect 5172 24216 5224 24225
rect 5356 24259 5408 24268
rect 5356 24225 5365 24259
rect 5365 24225 5399 24259
rect 5399 24225 5408 24259
rect 5356 24216 5408 24225
rect 7656 24259 7708 24268
rect 7656 24225 7665 24259
rect 7665 24225 7699 24259
rect 7699 24225 7708 24259
rect 7656 24216 7708 24225
rect 14464 24284 14516 24336
rect 15660 24284 15712 24336
rect 8484 24216 8536 24268
rect 10968 24259 11020 24268
rect 10968 24225 10977 24259
rect 10977 24225 11011 24259
rect 11011 24225 11020 24259
rect 10968 24216 11020 24225
rect 11428 24259 11480 24268
rect 11428 24225 11437 24259
rect 11437 24225 11471 24259
rect 11471 24225 11480 24259
rect 11428 24216 11480 24225
rect 2044 24148 2096 24200
rect 2964 24148 3016 24200
rect 7748 24148 7800 24200
rect 8760 24191 8812 24200
rect 4988 24080 5040 24132
rect 8760 24157 8769 24191
rect 8769 24157 8803 24191
rect 8803 24157 8812 24191
rect 8760 24148 8812 24157
rect 12256 24216 12308 24268
rect 13452 24259 13504 24268
rect 13452 24225 13461 24259
rect 13461 24225 13495 24259
rect 13495 24225 13504 24259
rect 13452 24216 13504 24225
rect 13544 24259 13596 24268
rect 13544 24225 13553 24259
rect 13553 24225 13587 24259
rect 13587 24225 13596 24259
rect 13544 24216 13596 24225
rect 16304 24216 16356 24268
rect 16764 24259 16816 24268
rect 16764 24225 16773 24259
rect 16773 24225 16807 24259
rect 16807 24225 16816 24259
rect 16764 24216 16816 24225
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 18880 24352 18932 24404
rect 22652 24352 22704 24404
rect 19156 24284 19208 24336
rect 12808 24191 12860 24200
rect 12808 24157 12817 24191
rect 12817 24157 12851 24191
rect 12851 24157 12860 24191
rect 12808 24148 12860 24157
rect 16672 24148 16724 24200
rect 18972 24216 19024 24268
rect 19340 24259 19392 24268
rect 19340 24225 19349 24259
rect 19349 24225 19383 24259
rect 19383 24225 19392 24259
rect 19340 24216 19392 24225
rect 21180 24259 21232 24268
rect 21180 24225 21189 24259
rect 21189 24225 21223 24259
rect 21223 24225 21232 24259
rect 21180 24216 21232 24225
rect 20352 24148 20404 24200
rect 21732 24148 21784 24200
rect 22928 24148 22980 24200
rect 9404 24080 9456 24132
rect 12900 24080 12952 24132
rect 18512 24080 18564 24132
rect 1860 24055 1912 24064
rect 1860 24021 1869 24055
rect 1869 24021 1903 24055
rect 1903 24021 1912 24055
rect 1860 24012 1912 24021
rect 3148 24012 3200 24064
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 12348 24012 12400 24064
rect 21456 24012 21508 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 1676 23851 1728 23860
rect 1676 23817 1685 23851
rect 1685 23817 1719 23851
rect 1719 23817 1728 23851
rect 1676 23808 1728 23817
rect 2044 23851 2096 23860
rect 2044 23817 2053 23851
rect 2053 23817 2087 23851
rect 2087 23817 2096 23851
rect 2044 23808 2096 23817
rect 5356 23808 5408 23860
rect 5908 23808 5960 23860
rect 6368 23851 6420 23860
rect 6368 23817 6377 23851
rect 6377 23817 6411 23851
rect 6411 23817 6420 23851
rect 6368 23808 6420 23817
rect 8484 23851 8536 23860
rect 8484 23817 8493 23851
rect 8493 23817 8527 23851
rect 8527 23817 8536 23851
rect 8484 23808 8536 23817
rect 9404 23808 9456 23860
rect 11428 23808 11480 23860
rect 11612 23808 11664 23860
rect 13544 23808 13596 23860
rect 16672 23808 16724 23860
rect 16764 23808 16816 23860
rect 4712 23740 4764 23792
rect 10968 23740 11020 23792
rect 12256 23740 12308 23792
rect 16120 23740 16172 23792
rect 16396 23740 16448 23792
rect 16948 23740 17000 23792
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 18880 23672 18932 23724
rect 20444 23808 20496 23860
rect 21180 23808 21232 23860
rect 22652 23851 22704 23860
rect 22652 23817 22661 23851
rect 22661 23817 22695 23851
rect 22695 23817 22704 23851
rect 22652 23808 22704 23817
rect 22928 23851 22980 23860
rect 22928 23817 22937 23851
rect 22937 23817 22971 23851
rect 22971 23817 22980 23851
rect 22928 23808 22980 23817
rect 2596 23604 2648 23656
rect 2964 23647 3016 23656
rect 2964 23613 2973 23647
rect 2973 23613 3007 23647
rect 3007 23613 3016 23647
rect 2964 23604 3016 23613
rect 3148 23647 3200 23656
rect 3148 23613 3157 23647
rect 3157 23613 3191 23647
rect 3191 23613 3200 23647
rect 3148 23604 3200 23613
rect 6368 23604 6420 23656
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 7748 23604 7800 23656
rect 8116 23647 8168 23656
rect 8116 23613 8125 23647
rect 8125 23613 8159 23647
rect 8159 23613 8168 23647
rect 8116 23604 8168 23613
rect 8760 23604 8812 23656
rect 12532 23604 12584 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 16120 23647 16172 23656
rect 16120 23613 16129 23647
rect 16129 23613 16163 23647
rect 16163 23613 16172 23647
rect 16120 23604 16172 23613
rect 2412 23536 2464 23588
rect 4620 23536 4672 23588
rect 12348 23536 12400 23588
rect 14648 23579 14700 23588
rect 14648 23545 14657 23579
rect 14657 23545 14691 23579
rect 14691 23545 14700 23579
rect 14648 23536 14700 23545
rect 16028 23536 16080 23588
rect 16764 23604 16816 23656
rect 19984 23672 20036 23724
rect 20168 23647 20220 23656
rect 20168 23613 20177 23647
rect 20177 23613 20211 23647
rect 20211 23613 20220 23647
rect 20352 23647 20404 23656
rect 20168 23604 20220 23613
rect 20352 23613 20361 23647
rect 20361 23613 20395 23647
rect 20395 23613 20404 23647
rect 20352 23604 20404 23613
rect 19156 23536 19208 23588
rect 21180 23579 21232 23588
rect 21180 23545 21189 23579
rect 21189 23545 21223 23579
rect 21223 23545 21232 23579
rect 21180 23536 21232 23545
rect 16212 23468 16264 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 2596 23307 2648 23316
rect 2596 23273 2605 23307
rect 2605 23273 2639 23307
rect 2639 23273 2648 23307
rect 2596 23264 2648 23273
rect 4436 23307 4488 23316
rect 4436 23273 4445 23307
rect 4445 23273 4479 23307
rect 4479 23273 4488 23307
rect 4436 23264 4488 23273
rect 5908 23264 5960 23316
rect 8116 23264 8168 23316
rect 11520 23264 11572 23316
rect 12256 23307 12308 23316
rect 4988 23239 5040 23248
rect 4988 23205 4997 23239
rect 4997 23205 5031 23239
rect 5031 23205 5040 23239
rect 4988 23196 5040 23205
rect 5724 23196 5776 23248
rect 6368 23196 6420 23248
rect 1584 23171 1636 23180
rect 1584 23137 1593 23171
rect 1593 23137 1627 23171
rect 1627 23137 1636 23171
rect 1584 23128 1636 23137
rect 1860 23128 1912 23180
rect 7196 23128 7248 23180
rect 8300 23128 8352 23180
rect 8576 23171 8628 23180
rect 8576 23137 8585 23171
rect 8585 23137 8619 23171
rect 8619 23137 8628 23171
rect 8576 23128 8628 23137
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 12256 23273 12265 23307
rect 12265 23273 12299 23307
rect 12299 23273 12308 23307
rect 12256 23264 12308 23273
rect 12808 23264 12860 23316
rect 16396 23264 16448 23316
rect 18512 23307 18564 23316
rect 18512 23273 18521 23307
rect 18521 23273 18555 23307
rect 18555 23273 18564 23307
rect 18512 23264 18564 23273
rect 19156 23307 19208 23316
rect 19156 23273 19165 23307
rect 19165 23273 19199 23307
rect 19199 23273 19208 23307
rect 19156 23264 19208 23273
rect 19984 23307 20036 23316
rect 19984 23273 19993 23307
rect 19993 23273 20027 23307
rect 20027 23273 20036 23307
rect 19984 23264 20036 23273
rect 16764 23196 16816 23248
rect 19340 23196 19392 23248
rect 20168 23196 20220 23248
rect 21180 23196 21232 23248
rect 2872 23060 2924 23112
rect 1676 22924 1728 22976
rect 2136 22924 2188 22976
rect 3608 22924 3660 22976
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 12624 23171 12676 23180
rect 12624 23137 12633 23171
rect 12633 23137 12667 23171
rect 12667 23137 12676 23171
rect 12624 23128 12676 23137
rect 13544 23128 13596 23180
rect 23020 23171 23072 23180
rect 23020 23137 23029 23171
rect 23029 23137 23063 23171
rect 23063 23137 23072 23171
rect 23020 23128 23072 23137
rect 13452 23103 13504 23112
rect 13452 23069 13461 23103
rect 13461 23069 13495 23103
rect 13495 23069 13504 23103
rect 13452 23060 13504 23069
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 16212 23103 16264 23112
rect 16212 23069 16221 23103
rect 16221 23069 16255 23103
rect 16255 23069 16264 23103
rect 16212 23060 16264 23069
rect 16580 23060 16632 23112
rect 22008 23060 22060 23112
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 11244 22992 11296 23044
rect 14648 22992 14700 23044
rect 21548 22992 21600 23044
rect 6092 22924 6144 22976
rect 8208 22924 8260 22976
rect 9956 22924 10008 22976
rect 10508 22924 10560 22976
rect 10968 22924 11020 22976
rect 15016 22924 15068 22976
rect 21180 22924 21232 22976
rect 22560 22924 22612 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 4988 22720 5040 22772
rect 5724 22763 5776 22772
rect 5724 22729 5733 22763
rect 5733 22729 5767 22763
rect 5767 22729 5776 22763
rect 5724 22720 5776 22729
rect 7196 22763 7248 22772
rect 7196 22729 7205 22763
rect 7205 22729 7239 22763
rect 7239 22729 7248 22763
rect 7196 22720 7248 22729
rect 10876 22720 10928 22772
rect 12440 22720 12492 22772
rect 16212 22720 16264 22772
rect 18512 22720 18564 22772
rect 23020 22763 23072 22772
rect 23020 22729 23029 22763
rect 23029 22729 23063 22763
rect 23063 22729 23072 22763
rect 23020 22720 23072 22729
rect 10508 22652 10560 22704
rect 13176 22695 13228 22704
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 10416 22584 10468 22636
rect 13176 22661 13185 22695
rect 13185 22661 13219 22695
rect 13219 22661 13228 22695
rect 13176 22652 13228 22661
rect 2136 22559 2188 22568
rect 2136 22525 2145 22559
rect 2145 22525 2179 22559
rect 2179 22525 2188 22559
rect 2136 22516 2188 22525
rect 8392 22559 8444 22568
rect 2872 22448 2924 22500
rect 4160 22491 4212 22500
rect 4160 22457 4169 22491
rect 4169 22457 4203 22491
rect 4203 22457 4212 22491
rect 4160 22448 4212 22457
rect 4620 22380 4672 22432
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 10968 22516 11020 22568
rect 11244 22559 11296 22568
rect 11244 22525 11253 22559
rect 11253 22525 11287 22559
rect 11287 22525 11296 22559
rect 11244 22516 11296 22525
rect 8484 22448 8536 22500
rect 10232 22491 10284 22500
rect 10232 22457 10241 22491
rect 10241 22457 10275 22491
rect 10275 22457 10284 22491
rect 10232 22448 10284 22457
rect 14924 22584 14976 22636
rect 15016 22584 15068 22636
rect 16028 22584 16080 22636
rect 20444 22627 20496 22636
rect 20444 22593 20453 22627
rect 20453 22593 20487 22627
rect 20487 22593 20496 22627
rect 20444 22584 20496 22593
rect 16304 22559 16356 22568
rect 16304 22525 16313 22559
rect 16313 22525 16347 22559
rect 16347 22525 16356 22559
rect 16304 22516 16356 22525
rect 17868 22516 17920 22568
rect 21180 22516 21232 22568
rect 21548 22559 21600 22568
rect 21548 22525 21557 22559
rect 21557 22525 21591 22559
rect 21591 22525 21600 22559
rect 21548 22516 21600 22525
rect 22008 22516 22060 22568
rect 14004 22448 14056 22500
rect 15292 22491 15344 22500
rect 15292 22457 15301 22491
rect 15301 22457 15335 22491
rect 15335 22457 15344 22491
rect 15292 22448 15344 22457
rect 6184 22380 6236 22432
rect 7932 22380 7984 22432
rect 8852 22380 8904 22432
rect 9956 22380 10008 22432
rect 10876 22380 10928 22432
rect 18052 22448 18104 22500
rect 19156 22448 19208 22500
rect 22836 22516 22888 22568
rect 21824 22380 21876 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 1584 22219 1636 22228
rect 1584 22185 1593 22219
rect 1593 22185 1627 22219
rect 1627 22185 1636 22219
rect 1584 22176 1636 22185
rect 2596 22040 2648 22092
rect 4160 22176 4212 22228
rect 7932 22176 7984 22228
rect 8576 22219 8628 22228
rect 8576 22185 8585 22219
rect 8585 22185 8619 22219
rect 8619 22185 8628 22219
rect 8576 22176 8628 22185
rect 11612 22219 11664 22228
rect 11612 22185 11621 22219
rect 11621 22185 11655 22219
rect 11655 22185 11664 22219
rect 11612 22176 11664 22185
rect 14004 22176 14056 22228
rect 5724 22108 5776 22160
rect 5356 22083 5408 22092
rect 5356 22049 5365 22083
rect 5365 22049 5399 22083
rect 5399 22049 5408 22083
rect 5356 22040 5408 22049
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8392 22040 8444 22092
rect 10232 22040 10284 22092
rect 10508 22083 10560 22092
rect 10508 22049 10517 22083
rect 10517 22049 10551 22083
rect 10551 22049 10560 22083
rect 10508 22040 10560 22049
rect 11244 22108 11296 22160
rect 12624 22108 12676 22160
rect 15292 22176 15344 22228
rect 16764 22219 16816 22228
rect 16764 22185 16773 22219
rect 16773 22185 16807 22219
rect 16807 22185 16816 22219
rect 16764 22176 16816 22185
rect 18604 22108 18656 22160
rect 19984 22108 20036 22160
rect 22100 22108 22152 22160
rect 10968 22040 11020 22092
rect 12992 22040 13044 22092
rect 14188 22083 14240 22092
rect 14188 22049 14197 22083
rect 14197 22049 14231 22083
rect 14231 22049 14240 22083
rect 14188 22040 14240 22049
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 17868 22083 17920 22092
rect 2320 21972 2372 22024
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 12624 21972 12676 22024
rect 13176 21972 13228 22024
rect 14740 21972 14792 22024
rect 15936 21972 15988 22024
rect 17868 22049 17877 22083
rect 17877 22049 17911 22083
rect 17911 22049 17920 22083
rect 17868 22040 17920 22049
rect 21180 22083 21232 22092
rect 21180 22049 21189 22083
rect 21189 22049 21223 22083
rect 21223 22049 21232 22083
rect 21180 22040 21232 22049
rect 21548 22040 21600 22092
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 18144 21972 18196 21981
rect 9680 21904 9732 21956
rect 2504 21836 2556 21888
rect 22192 21836 22244 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 2872 21632 2924 21684
rect 5356 21632 5408 21684
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 11980 21675 12032 21684
rect 11980 21641 11989 21675
rect 11989 21641 12023 21675
rect 12023 21641 12032 21675
rect 11980 21632 12032 21641
rect 16304 21632 16356 21684
rect 18144 21632 18196 21684
rect 22836 21632 22888 21684
rect 5632 21564 5684 21616
rect 6092 21564 6144 21616
rect 2504 21496 2556 21548
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 10416 21496 10468 21548
rect 18604 21564 18656 21616
rect 12992 21496 13044 21548
rect 2136 21428 2188 21480
rect 2596 21471 2648 21480
rect 2596 21437 2605 21471
rect 2605 21437 2639 21471
rect 2639 21437 2648 21471
rect 2596 21428 2648 21437
rect 2320 21360 2372 21412
rect 2228 21335 2280 21344
rect 2228 21301 2237 21335
rect 2237 21301 2271 21335
rect 2271 21301 2280 21335
rect 2228 21292 2280 21301
rect 8576 21428 8628 21480
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 18328 21428 18380 21480
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 10140 21360 10192 21412
rect 13360 21360 13412 21412
rect 16948 21360 17000 21412
rect 18604 21360 18656 21412
rect 21548 21539 21600 21548
rect 21548 21505 21557 21539
rect 21557 21505 21591 21539
rect 21591 21505 21600 21539
rect 21548 21496 21600 21505
rect 23020 21496 23072 21548
rect 19248 21471 19300 21480
rect 19248 21437 19257 21471
rect 19257 21437 19291 21471
rect 19291 21437 19300 21471
rect 19248 21428 19300 21437
rect 22192 21471 22244 21480
rect 4620 21292 4672 21344
rect 14924 21335 14976 21344
rect 14924 21301 14933 21335
rect 14933 21301 14967 21335
rect 14967 21301 14976 21335
rect 16580 21335 16632 21344
rect 14924 21292 14976 21301
rect 16580 21301 16589 21335
rect 16589 21301 16623 21335
rect 16623 21301 16632 21335
rect 16580 21292 16632 21301
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 22836 21428 22888 21480
rect 21088 21292 21140 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 3608 21131 3660 21140
rect 3608 21097 3617 21131
rect 3617 21097 3651 21131
rect 3651 21097 3660 21131
rect 3608 21088 3660 21097
rect 7840 21088 7892 21140
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 8852 21131 8904 21140
rect 8852 21097 8861 21131
rect 8861 21097 8895 21131
rect 8895 21097 8904 21131
rect 8852 21088 8904 21097
rect 12348 21131 12400 21140
rect 12348 21097 12357 21131
rect 12357 21097 12391 21131
rect 12391 21097 12400 21131
rect 12348 21088 12400 21097
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 18328 21131 18380 21140
rect 18328 21097 18337 21131
rect 18337 21097 18371 21131
rect 18371 21097 18380 21131
rect 18328 21088 18380 21097
rect 21180 21088 21232 21140
rect 22008 21088 22060 21140
rect 22560 21088 22612 21140
rect 1676 21020 1728 21072
rect 5724 21020 5776 21072
rect 6092 21020 6144 21072
rect 7656 21020 7708 21072
rect 10508 21020 10560 21072
rect 12992 21020 13044 21072
rect 18144 21020 18196 21072
rect 21824 21063 21876 21072
rect 21824 21029 21833 21063
rect 21833 21029 21867 21063
rect 21867 21029 21876 21063
rect 21824 21020 21876 21029
rect 22376 21020 22428 21072
rect 2228 20952 2280 21004
rect 2320 20995 2372 21004
rect 2320 20961 2329 20995
rect 2329 20961 2363 20995
rect 2363 20961 2372 20995
rect 2504 20995 2556 21004
rect 2320 20952 2372 20961
rect 2504 20961 2513 20995
rect 2513 20961 2547 20995
rect 2547 20961 2556 20995
rect 2504 20952 2556 20961
rect 4620 20952 4672 21004
rect 10416 20995 10468 21004
rect 10416 20961 10425 20995
rect 10425 20961 10459 20995
rect 10459 20961 10468 20995
rect 10416 20952 10468 20961
rect 11428 20952 11480 21004
rect 13820 20952 13872 21004
rect 14188 20995 14240 21004
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 14924 20952 14976 21004
rect 16488 20995 16540 21004
rect 16488 20961 16497 20995
rect 16497 20961 16531 20995
rect 16531 20961 16540 20995
rect 16488 20952 16540 20961
rect 16948 20995 17000 21004
rect 16948 20961 16957 20995
rect 16957 20961 16991 20995
rect 16991 20961 17000 20995
rect 16948 20952 17000 20961
rect 18880 20952 18932 21004
rect 20444 20952 20496 21004
rect 1676 20927 1728 20936
rect 1676 20893 1685 20927
rect 1685 20893 1719 20927
rect 1719 20893 1728 20927
rect 1676 20884 1728 20893
rect 2412 20816 2464 20868
rect 3516 20816 3568 20868
rect 2044 20748 2096 20800
rect 3608 20748 3660 20800
rect 6092 20884 6144 20936
rect 17776 20884 17828 20936
rect 19248 20884 19300 20936
rect 8576 20816 8628 20868
rect 14740 20816 14792 20868
rect 19616 20816 19668 20868
rect 21456 20884 21508 20936
rect 23020 20884 23072 20936
rect 18604 20791 18656 20800
rect 18604 20757 18613 20791
rect 18613 20757 18647 20791
rect 18647 20757 18656 20791
rect 18604 20748 18656 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 2136 20544 2188 20596
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 5724 20544 5776 20596
rect 10140 20544 10192 20596
rect 16488 20544 16540 20596
rect 16948 20544 17000 20596
rect 18880 20544 18932 20596
rect 21824 20544 21876 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 10416 20476 10468 20528
rect 8484 20408 8536 20460
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 14648 20408 14700 20460
rect 16304 20408 16356 20460
rect 20352 20408 20404 20460
rect 20444 20408 20496 20460
rect 2044 20340 2096 20392
rect 3516 20340 3568 20392
rect 6092 20340 6144 20392
rect 7840 20383 7892 20392
rect 7840 20349 7849 20383
rect 7849 20349 7883 20383
rect 7883 20349 7892 20383
rect 7840 20340 7892 20349
rect 8576 20272 8628 20324
rect 9864 20315 9916 20324
rect 9864 20281 9873 20315
rect 9873 20281 9907 20315
rect 9907 20281 9916 20315
rect 9864 20272 9916 20281
rect 4620 20204 4672 20256
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 13728 20340 13780 20392
rect 19616 20383 19668 20392
rect 19616 20349 19625 20383
rect 19625 20349 19659 20383
rect 19659 20349 19668 20383
rect 19616 20340 19668 20349
rect 14280 20315 14332 20324
rect 14280 20281 14289 20315
rect 14289 20281 14323 20315
rect 14323 20281 14332 20315
rect 14280 20272 14332 20281
rect 14740 20272 14792 20324
rect 11428 20204 11480 20256
rect 12992 20204 13044 20256
rect 13728 20204 13780 20256
rect 13820 20204 13872 20256
rect 14464 20204 14516 20256
rect 20352 20272 20404 20324
rect 22100 20204 22152 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 3516 20000 3568 20052
rect 14740 20000 14792 20052
rect 16488 20000 16540 20052
rect 2412 19975 2464 19984
rect 2412 19941 2421 19975
rect 2421 19941 2455 19975
rect 2455 19941 2464 19975
rect 2412 19932 2464 19941
rect 6828 19932 6880 19984
rect 2136 19864 2188 19916
rect 4068 19864 4120 19916
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 9312 19864 9364 19916
rect 9864 19864 9916 19916
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 12992 19864 13044 19916
rect 15936 19864 15988 19916
rect 20352 20000 20404 20052
rect 16948 19932 17000 19984
rect 16764 19864 16816 19916
rect 20444 19932 20496 19984
rect 22560 19975 22612 19984
rect 22560 19941 22569 19975
rect 22569 19941 22603 19975
rect 22603 19941 22612 19975
rect 22560 19932 22612 19941
rect 17776 19907 17828 19916
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 17960 19907 18012 19916
rect 17960 19873 17969 19907
rect 17969 19873 18003 19907
rect 18003 19873 18012 19907
rect 17960 19864 18012 19873
rect 5724 19796 5776 19848
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 8116 19839 8168 19848
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 11152 19796 11204 19848
rect 16028 19839 16080 19848
rect 15292 19728 15344 19780
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 18328 19864 18380 19916
rect 19432 19864 19484 19916
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 22192 19864 22244 19916
rect 22744 19864 22796 19916
rect 18604 19796 18656 19848
rect 16120 19728 16172 19780
rect 3516 19703 3568 19712
rect 3516 19669 3525 19703
rect 3525 19669 3559 19703
rect 3559 19669 3568 19703
rect 3516 19660 3568 19669
rect 9312 19703 9364 19712
rect 9312 19669 9321 19703
rect 9321 19669 9355 19703
rect 9355 19669 9364 19703
rect 9312 19660 9364 19669
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 12072 19660 12124 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 18512 19660 18564 19712
rect 21456 19660 21508 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 3516 19456 3568 19508
rect 5356 19456 5408 19508
rect 6368 19456 6420 19508
rect 7840 19456 7892 19508
rect 8576 19456 8628 19508
rect 16764 19499 16816 19508
rect 16764 19465 16773 19499
rect 16773 19465 16807 19499
rect 16807 19465 16816 19499
rect 16764 19456 16816 19465
rect 19064 19456 19116 19508
rect 21088 19456 21140 19508
rect 22376 19456 22428 19508
rect 22744 19499 22796 19508
rect 22744 19465 22753 19499
rect 22753 19465 22787 19499
rect 22787 19465 22796 19499
rect 22744 19456 22796 19465
rect 9864 19320 9916 19372
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 2228 19252 2280 19304
rect 3516 19252 3568 19304
rect 5724 19295 5776 19304
rect 2412 19116 2464 19168
rect 4068 19184 4120 19236
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 6276 19252 6328 19304
rect 7104 19252 7156 19304
rect 8116 19252 8168 19304
rect 11520 19320 11572 19372
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 19524 19320 19576 19372
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 11152 19295 11204 19304
rect 10324 19184 10376 19236
rect 11152 19261 11161 19295
rect 11161 19261 11195 19295
rect 11195 19261 11204 19295
rect 11152 19252 11204 19261
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 12900 19252 12952 19261
rect 14004 19252 14056 19304
rect 14464 19252 14516 19304
rect 11520 19227 11572 19236
rect 11520 19193 11529 19227
rect 11529 19193 11563 19227
rect 11563 19193 11572 19227
rect 11520 19184 11572 19193
rect 12716 19184 12768 19236
rect 14280 19184 14332 19236
rect 16028 19252 16080 19304
rect 16580 19295 16632 19304
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 21088 19252 21140 19304
rect 22284 19252 22336 19304
rect 17316 19184 17368 19236
rect 19248 19184 19300 19236
rect 11428 19116 11480 19168
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 16028 19159 16080 19168
rect 16028 19125 16037 19159
rect 16037 19125 16071 19159
rect 16071 19125 16080 19159
rect 16028 19116 16080 19125
rect 16120 19116 16172 19168
rect 21732 19116 21784 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 2320 18912 2372 18964
rect 5724 18912 5776 18964
rect 6368 18912 6420 18964
rect 6828 18912 6880 18964
rect 9312 18955 9364 18964
rect 9312 18921 9321 18955
rect 9321 18921 9355 18955
rect 9355 18921 9364 18955
rect 9312 18912 9364 18921
rect 10508 18912 10560 18964
rect 11152 18912 11204 18964
rect 14096 18912 14148 18964
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 17776 18912 17828 18964
rect 19248 18955 19300 18964
rect 19248 18921 19257 18955
rect 19257 18921 19291 18955
rect 19291 18921 19300 18955
rect 19248 18912 19300 18921
rect 19432 18912 19484 18964
rect 2136 18844 2188 18896
rect 5356 18844 5408 18896
rect 1676 18776 1728 18828
rect 3056 18776 3108 18828
rect 5080 18776 5132 18828
rect 7104 18887 7156 18896
rect 7104 18853 7113 18887
rect 7113 18853 7147 18887
rect 7147 18853 7156 18887
rect 7104 18844 7156 18853
rect 12716 18887 12768 18896
rect 12716 18853 12725 18887
rect 12725 18853 12759 18887
rect 12759 18853 12768 18887
rect 12716 18844 12768 18853
rect 17960 18844 18012 18896
rect 21824 18844 21876 18896
rect 22744 18844 22796 18896
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 5632 18708 5684 18760
rect 4620 18640 4672 18692
rect 7840 18776 7892 18828
rect 12072 18776 12124 18828
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 19064 18819 19116 18828
rect 19064 18785 19073 18819
rect 19073 18785 19107 18819
rect 19107 18785 19116 18819
rect 19064 18776 19116 18785
rect 10968 18751 11020 18760
rect 3148 18615 3200 18624
rect 3148 18581 3157 18615
rect 3157 18581 3191 18615
rect 3191 18581 3200 18615
rect 3148 18572 3200 18581
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 16396 18708 16448 18760
rect 20444 18708 20496 18760
rect 21364 18751 21416 18760
rect 11060 18572 11112 18624
rect 11428 18572 11480 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 14004 18572 14056 18624
rect 18236 18572 18288 18624
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 21456 18572 21508 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 5080 18411 5132 18420
rect 5080 18377 5089 18411
rect 5089 18377 5123 18411
rect 5123 18377 5132 18411
rect 5080 18368 5132 18377
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 5816 18368 5868 18420
rect 10324 18368 10376 18420
rect 21364 18368 21416 18420
rect 4804 18300 4856 18352
rect 6276 18300 6328 18352
rect 10968 18343 11020 18352
rect 10968 18309 10977 18343
rect 10977 18309 11011 18343
rect 11011 18309 11020 18343
rect 10968 18300 11020 18309
rect 19432 18300 19484 18352
rect 2044 18232 2096 18284
rect 4068 18232 4120 18284
rect 2596 18096 2648 18148
rect 2964 18096 3016 18148
rect 5356 18232 5408 18284
rect 8760 18232 8812 18284
rect 7840 18207 7892 18216
rect 7840 18173 7849 18207
rect 7849 18173 7883 18207
rect 7883 18173 7892 18207
rect 9864 18207 9916 18216
rect 7840 18164 7892 18173
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 14096 18232 14148 18284
rect 15108 18232 15160 18284
rect 15936 18232 15988 18284
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 10324 18096 10376 18148
rect 14740 18139 14792 18148
rect 14740 18105 14749 18139
rect 14749 18105 14783 18139
rect 14783 18105 14792 18139
rect 14740 18096 14792 18105
rect 15752 18096 15804 18148
rect 8024 18071 8076 18080
rect 8024 18037 8033 18071
rect 8033 18037 8067 18071
rect 8067 18037 8076 18071
rect 8024 18028 8076 18037
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 13084 18028 13136 18080
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 19064 18071 19116 18080
rect 19064 18037 19073 18071
rect 19073 18037 19107 18071
rect 19107 18037 19116 18071
rect 19064 18028 19116 18037
rect 22468 18071 22520 18080
rect 22468 18037 22477 18071
rect 22477 18037 22511 18071
rect 22511 18037 22520 18071
rect 22468 18028 22520 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 2964 17824 3016 17876
rect 8300 17824 8352 17876
rect 10048 17824 10100 17876
rect 12072 17824 12124 17876
rect 15752 17824 15804 17876
rect 19156 17824 19208 17876
rect 19432 17824 19484 17876
rect 20904 17824 20956 17876
rect 2044 17756 2096 17808
rect 3056 17799 3108 17808
rect 3056 17765 3065 17799
rect 3065 17765 3099 17799
rect 3099 17765 3108 17799
rect 3056 17756 3108 17765
rect 13084 17799 13136 17808
rect 13084 17765 13093 17799
rect 13093 17765 13127 17799
rect 13127 17765 13136 17799
rect 13084 17756 13136 17765
rect 14924 17799 14976 17808
rect 14924 17765 14933 17799
rect 14933 17765 14967 17799
rect 14967 17765 14976 17799
rect 14924 17756 14976 17765
rect 22468 17756 22520 17808
rect 3240 17688 3292 17740
rect 4620 17688 4672 17740
rect 5356 17620 5408 17672
rect 6828 17688 6880 17740
rect 6920 17688 6972 17740
rect 8208 17688 8260 17740
rect 8576 17688 8628 17740
rect 9036 17688 9088 17740
rect 11428 17688 11480 17740
rect 11704 17688 11756 17740
rect 13268 17688 13320 17740
rect 16488 17731 16540 17740
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 12072 17620 12124 17672
rect 14004 17620 14056 17672
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16488 17697 16497 17731
rect 16497 17697 16531 17731
rect 16531 17697 16540 17731
rect 16488 17688 16540 17697
rect 17316 17688 17368 17740
rect 17776 17688 17828 17740
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 18972 17620 19024 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 21732 17663 21784 17672
rect 21732 17629 21741 17663
rect 21741 17629 21775 17663
rect 21775 17629 21784 17663
rect 21732 17620 21784 17629
rect 22376 17620 22428 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 4988 17484 5040 17536
rect 9312 17484 9364 17536
rect 9864 17484 9916 17536
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 11060 17484 11112 17493
rect 11520 17484 11572 17536
rect 17500 17484 17552 17536
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 20996 17484 21048 17536
rect 21824 17484 21876 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 5448 17280 5500 17332
rect 6920 17280 6972 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 15936 17280 15988 17332
rect 16488 17323 16540 17332
rect 16488 17289 16497 17323
rect 16497 17289 16531 17323
rect 16531 17289 16540 17323
rect 16488 17280 16540 17289
rect 17316 17323 17368 17332
rect 17316 17289 17325 17323
rect 17325 17289 17359 17323
rect 17359 17289 17368 17323
rect 17316 17280 17368 17289
rect 22468 17280 22520 17332
rect 14464 17212 14516 17264
rect 14740 17212 14792 17264
rect 21732 17212 21784 17264
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 12900 17144 12952 17196
rect 18604 17144 18656 17196
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 2044 17076 2096 17128
rect 4068 17076 4120 17128
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 6644 17076 6696 17128
rect 9312 17076 9364 17128
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 13176 17076 13228 17128
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 14096 17119 14148 17128
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 3148 17008 3200 17060
rect 3700 17008 3752 17060
rect 6092 17008 6144 17060
rect 10784 17008 10836 17060
rect 14924 17076 14976 17128
rect 17500 17076 17552 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 21088 17119 21140 17128
rect 21088 17085 21097 17119
rect 21097 17085 21131 17119
rect 21131 17085 21140 17119
rect 21088 17076 21140 17085
rect 21180 17076 21232 17128
rect 22652 17076 22704 17128
rect 14832 17008 14884 17060
rect 16396 17008 16448 17060
rect 18972 17008 19024 17060
rect 20260 17051 20312 17060
rect 20260 17017 20269 17051
rect 20269 17017 20303 17051
rect 20303 17017 20312 17051
rect 20260 17008 20312 17017
rect 4620 16940 4672 16992
rect 5080 16940 5132 16992
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 10232 16940 10284 16992
rect 11428 16940 11480 16992
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 21456 16940 21508 16992
rect 22928 16983 22980 16992
rect 22928 16949 22937 16983
rect 22937 16949 22971 16983
rect 22971 16949 22980 16983
rect 22928 16940 22980 16949
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 3148 16736 3200 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3700 16779 3752 16788
rect 3240 16736 3292 16745
rect 3700 16745 3709 16779
rect 3709 16745 3743 16779
rect 3743 16745 3752 16779
rect 3700 16736 3752 16745
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 8024 16736 8076 16788
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 14004 16736 14056 16788
rect 14096 16736 14148 16788
rect 14832 16779 14884 16788
rect 14832 16745 14841 16779
rect 14841 16745 14875 16779
rect 14875 16745 14884 16779
rect 14832 16736 14884 16745
rect 1676 16668 1728 16720
rect 2320 16668 2372 16720
rect 10784 16668 10836 16720
rect 11520 16668 11572 16720
rect 4988 16600 5040 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5908 16643 5960 16652
rect 5448 16600 5500 16609
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 5908 16600 5960 16609
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 8576 16643 8628 16652
rect 8576 16609 8585 16643
rect 8585 16609 8619 16643
rect 8619 16609 8628 16643
rect 9864 16643 9916 16652
rect 8576 16600 8628 16609
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 2504 16532 2556 16584
rect 4896 16464 4948 16516
rect 1676 16396 1728 16448
rect 4068 16396 4120 16448
rect 8760 16439 8812 16448
rect 8760 16405 8769 16439
rect 8769 16405 8803 16439
rect 8803 16405 8812 16439
rect 8760 16396 8812 16405
rect 10232 16396 10284 16448
rect 15108 16600 15160 16652
rect 18236 16736 18288 16788
rect 18972 16736 19024 16788
rect 16488 16668 16540 16720
rect 17500 16711 17552 16720
rect 17500 16677 17509 16711
rect 17509 16677 17543 16711
rect 17543 16677 17552 16711
rect 17500 16668 17552 16677
rect 20444 16668 20496 16720
rect 21088 16668 21140 16720
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 19432 16600 19484 16652
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 11060 16532 11112 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 22376 16575 22428 16584
rect 22376 16541 22385 16575
rect 22385 16541 22419 16575
rect 22419 16541 22428 16575
rect 22376 16532 22428 16541
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 18788 16464 18840 16516
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 20536 16439 20588 16448
rect 20536 16405 20545 16439
rect 20545 16405 20579 16439
rect 20579 16405 20588 16439
rect 20536 16396 20588 16405
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 6092 16192 6144 16244
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 11520 16192 11572 16244
rect 12900 16192 12952 16244
rect 15108 16235 15160 16244
rect 15108 16201 15117 16235
rect 15117 16201 15151 16235
rect 15151 16201 15160 16235
rect 15108 16192 15160 16201
rect 16488 16235 16540 16244
rect 16488 16201 16497 16235
rect 16497 16201 16531 16235
rect 16531 16201 16540 16235
rect 16488 16192 16540 16201
rect 17776 16192 17828 16244
rect 20536 16192 20588 16244
rect 22652 16192 22704 16244
rect 21180 16124 21232 16176
rect 22560 16124 22612 16176
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 5356 16031 5408 16040
rect 2596 15920 2648 15972
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 5908 16056 5960 16108
rect 7472 16099 7524 16108
rect 7472 16065 7481 16099
rect 7481 16065 7515 16099
rect 7515 16065 7524 16099
rect 7472 16056 7524 16065
rect 8484 16056 8536 16108
rect 11152 16056 11204 16108
rect 15752 16056 15804 16108
rect 19248 16056 19300 16108
rect 22376 16056 22428 16108
rect 6092 15988 6144 16040
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 10140 15988 10192 16040
rect 6644 15920 6696 15972
rect 8024 15920 8076 15972
rect 10416 15920 10468 15972
rect 13176 15988 13228 16040
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 22284 15988 22336 16040
rect 11060 15852 11112 15904
rect 14188 15852 14240 15904
rect 18788 15920 18840 15972
rect 17868 15852 17920 15904
rect 20904 15920 20956 15972
rect 23388 15852 23440 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 7472 15648 7524 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 12532 15648 12584 15700
rect 20996 15648 21048 15700
rect 1860 15512 1912 15564
rect 2228 15512 2280 15564
rect 2596 15580 2648 15632
rect 4896 15623 4948 15632
rect 4896 15589 4905 15623
rect 4905 15589 4939 15623
rect 4939 15589 4948 15623
rect 4896 15580 4948 15589
rect 5540 15580 5592 15632
rect 6644 15623 6696 15632
rect 6644 15589 6653 15623
rect 6653 15589 6687 15623
rect 6687 15589 6696 15623
rect 6644 15580 6696 15589
rect 17040 15580 17092 15632
rect 20260 15580 20312 15632
rect 22560 15623 22612 15632
rect 22560 15589 22569 15623
rect 22569 15589 22603 15623
rect 22603 15589 22612 15623
rect 22560 15580 22612 15589
rect 2504 15555 2556 15564
rect 2504 15521 2513 15555
rect 2513 15521 2547 15555
rect 2547 15521 2556 15555
rect 2504 15512 2556 15521
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 20628 15512 20680 15564
rect 21916 15512 21968 15564
rect 22376 15512 22428 15564
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 6276 15444 6328 15496
rect 7012 15444 7064 15496
rect 7196 15444 7248 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 2504 15376 2556 15428
rect 14832 15376 14884 15428
rect 1676 15308 1728 15360
rect 5448 15308 5500 15360
rect 10600 15308 10652 15360
rect 13544 15308 13596 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 18512 15308 18564 15360
rect 19432 15308 19484 15360
rect 19892 15308 19944 15360
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 4896 15104 4948 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 15844 15104 15896 15156
rect 18420 15104 18472 15156
rect 20628 15104 20680 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 22376 15104 22428 15156
rect 3608 15036 3660 15088
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 2044 14900 2096 14952
rect 3608 14900 3660 14952
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 5632 14900 5684 14952
rect 4344 14832 4396 14884
rect 7840 14832 7892 14884
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 8576 14943 8628 14952
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 12808 14900 12860 14952
rect 13360 14900 13412 14952
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 18420 14943 18472 14952
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 18512 14900 18564 14952
rect 20904 14943 20956 14952
rect 20904 14909 20913 14943
rect 20913 14909 20947 14943
rect 20947 14909 20956 14943
rect 20904 14900 20956 14909
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 16396 14875 16448 14884
rect 16396 14841 16405 14875
rect 16405 14841 16439 14875
rect 16439 14841 16448 14875
rect 16396 14832 16448 14841
rect 19248 14832 19300 14884
rect 20260 14832 20312 14884
rect 8760 14764 8812 14816
rect 10048 14764 10100 14816
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 15936 14807 15988 14816
rect 15936 14773 15945 14807
rect 15945 14773 15979 14807
rect 15979 14773 15988 14807
rect 15936 14764 15988 14773
rect 22192 14764 22244 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 3608 14560 3660 14612
rect 5632 14603 5684 14612
rect 5632 14569 5641 14603
rect 5641 14569 5675 14603
rect 5675 14569 5684 14603
rect 5632 14560 5684 14569
rect 8484 14603 8536 14612
rect 8484 14569 8493 14603
rect 8493 14569 8527 14603
rect 8527 14569 8536 14603
rect 8484 14560 8536 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 14464 14560 14516 14612
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 11796 14492 11848 14544
rect 14924 14535 14976 14544
rect 14924 14501 14933 14535
rect 14933 14501 14967 14535
rect 14967 14501 14976 14535
rect 14924 14492 14976 14501
rect 15108 14492 15160 14544
rect 18788 14560 18840 14612
rect 4344 14424 4396 14476
rect 4988 14424 5040 14476
rect 7472 14424 7524 14476
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 9680 14424 9732 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 10692 14424 10744 14476
rect 14188 14467 14240 14476
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 19156 14492 19208 14544
rect 2412 14356 2464 14408
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 7748 14356 7800 14408
rect 11060 14399 11112 14408
rect 2780 14288 2832 14340
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 8024 14288 8076 14340
rect 9864 14288 9916 14340
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 7196 14220 7248 14229
rect 10232 14263 10284 14272
rect 10232 14229 10241 14263
rect 10241 14229 10275 14263
rect 10275 14229 10284 14263
rect 10232 14220 10284 14229
rect 18512 14424 18564 14476
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 19340 14467 19392 14476
rect 19340 14433 19349 14467
rect 19349 14433 19383 14467
rect 19383 14433 19392 14467
rect 19340 14424 19392 14433
rect 22192 14492 22244 14544
rect 23388 14535 23440 14544
rect 23388 14501 23397 14535
rect 23397 14501 23431 14535
rect 23431 14501 23440 14535
rect 23388 14492 23440 14501
rect 20260 14424 20312 14476
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 16120 14356 16172 14408
rect 18420 14356 18472 14408
rect 18880 14356 18932 14408
rect 21364 14399 21416 14408
rect 21364 14365 21373 14399
rect 21373 14365 21407 14399
rect 21407 14365 21416 14399
rect 21364 14356 21416 14365
rect 22100 14356 22152 14408
rect 17224 14220 17276 14272
rect 19984 14220 20036 14272
rect 20904 14220 20956 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 1676 14016 1728 14068
rect 4988 14059 5040 14068
rect 4988 14025 4997 14059
rect 4997 14025 5031 14059
rect 5031 14025 5040 14059
rect 4988 14016 5040 14025
rect 7472 14016 7524 14068
rect 2044 13880 2096 13932
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 6276 13880 6328 13932
rect 6920 13880 6972 13932
rect 7380 13880 7432 13932
rect 7748 13880 7800 13932
rect 2136 13812 2188 13864
rect 4068 13812 4120 13864
rect 5632 13812 5684 13864
rect 9220 13812 9272 13864
rect 10232 14016 10284 14068
rect 11796 14016 11848 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 18420 14016 18472 14068
rect 22192 14016 22244 14068
rect 10692 13991 10744 14000
rect 10692 13957 10701 13991
rect 10701 13957 10735 13991
rect 10735 13957 10744 13991
rect 10692 13948 10744 13957
rect 11336 13948 11388 14000
rect 15844 13948 15896 14000
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 11888 13880 11940 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 12716 13812 12768 13864
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 13360 13855 13412 13864
rect 12900 13812 12952 13821
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 13544 13855 13596 13864
rect 13544 13821 13553 13855
rect 13553 13821 13587 13855
rect 13587 13821 13596 13855
rect 13544 13812 13596 13821
rect 2964 13787 3016 13796
rect 2964 13753 2973 13787
rect 2973 13753 3007 13787
rect 3007 13753 3016 13787
rect 2964 13744 3016 13753
rect 4712 13787 4764 13796
rect 4712 13753 4721 13787
rect 4721 13753 4755 13787
rect 4755 13753 4764 13787
rect 4712 13744 4764 13753
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 7932 13744 7984 13796
rect 16396 13812 16448 13864
rect 16672 13880 16724 13932
rect 19432 13948 19484 14000
rect 20904 13948 20956 14000
rect 21364 13948 21416 14000
rect 22928 13948 22980 14000
rect 19984 13880 20036 13932
rect 19156 13812 19208 13864
rect 20076 13855 20128 13864
rect 16948 13744 17000 13796
rect 18788 13744 18840 13796
rect 19248 13744 19300 13796
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 15200 13719 15252 13728
rect 15200 13685 15209 13719
rect 15209 13685 15243 13719
rect 15243 13685 15252 13719
rect 15200 13676 15252 13685
rect 15568 13719 15620 13728
rect 15568 13685 15577 13719
rect 15577 13685 15611 13719
rect 15611 13685 15620 13719
rect 15568 13676 15620 13685
rect 19340 13676 19392 13728
rect 20076 13676 20128 13728
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 2596 13515 2648 13524
rect 2596 13481 2605 13515
rect 2605 13481 2639 13515
rect 2639 13481 2648 13515
rect 2596 13472 2648 13481
rect 2964 13472 3016 13524
rect 4068 13404 4120 13456
rect 7288 13472 7340 13524
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 13360 13472 13412 13524
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 15200 13472 15252 13524
rect 15752 13472 15804 13524
rect 16948 13472 17000 13524
rect 19156 13515 19208 13524
rect 19156 13481 19165 13515
rect 19165 13481 19199 13515
rect 19199 13481 19208 13515
rect 19156 13472 19208 13481
rect 19340 13472 19392 13524
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 7656 13404 7708 13456
rect 7932 13404 7984 13456
rect 9772 13404 9824 13456
rect 10600 13404 10652 13456
rect 11888 13447 11940 13456
rect 11888 13413 11897 13447
rect 11897 13413 11931 13447
rect 11931 13413 11940 13447
rect 11888 13404 11940 13413
rect 12716 13404 12768 13456
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7196 13336 7248 13388
rect 7472 13336 7524 13388
rect 7748 13336 7800 13388
rect 8024 13379 8076 13388
rect 8024 13345 8033 13379
rect 8033 13345 8067 13379
rect 8067 13345 8076 13379
rect 8024 13336 8076 13345
rect 15568 13336 15620 13388
rect 15844 13336 15896 13388
rect 19248 13404 19300 13456
rect 21364 13404 21416 13456
rect 16764 13336 16816 13388
rect 17868 13336 17920 13388
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 22100 13404 22152 13456
rect 5172 13200 5224 13252
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 15660 13200 15712 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 2136 13132 2188 13184
rect 3608 13132 3660 13184
rect 7564 13132 7616 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 18972 13132 19024 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 2688 12928 2740 12980
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 4620 12928 4672 12980
rect 5172 12928 5224 12980
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 7104 12928 7156 12980
rect 8208 12928 8260 12980
rect 10600 12928 10652 12980
rect 15844 12928 15896 12980
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 4712 12860 4764 12912
rect 7472 12860 7524 12912
rect 8024 12792 8076 12844
rect 19248 12792 19300 12844
rect 5356 12767 5408 12776
rect 1676 12724 1728 12733
rect 3608 12656 3660 12708
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 14372 12767 14424 12776
rect 14372 12733 14381 12767
rect 14381 12733 14415 12767
rect 14415 12733 14424 12767
rect 14372 12724 14424 12733
rect 14464 12724 14516 12776
rect 15568 12724 15620 12776
rect 16304 12724 16356 12776
rect 17224 12724 17276 12776
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 21456 12724 21508 12776
rect 22468 12724 22520 12776
rect 23388 12724 23440 12776
rect 6920 12656 6972 12708
rect 9864 12656 9916 12708
rect 2780 12588 2832 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 10600 12588 10652 12640
rect 12624 12656 12676 12708
rect 14924 12656 14976 12708
rect 15476 12656 15528 12708
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 18972 12656 19024 12708
rect 22008 12699 22060 12708
rect 22008 12665 22017 12699
rect 22017 12665 22051 12699
rect 22051 12665 22060 12699
rect 22008 12656 22060 12665
rect 21548 12588 21600 12640
rect 21732 12588 21784 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 2596 12384 2648 12436
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 8208 12427 8260 12436
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 9772 12384 9824 12436
rect 12624 12427 12676 12436
rect 1124 12248 1176 12300
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 5080 12248 5132 12300
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 16304 12427 16356 12436
rect 16304 12393 16313 12427
rect 16313 12393 16347 12427
rect 16347 12393 16356 12427
rect 16304 12384 16356 12393
rect 17224 12384 17276 12436
rect 18880 12384 18932 12436
rect 21732 12316 21784 12368
rect 22100 12316 22152 12368
rect 23388 12359 23440 12368
rect 23388 12325 23397 12359
rect 23397 12325 23431 12359
rect 23431 12325 23440 12359
rect 23388 12316 23440 12325
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 1492 12180 1544 12232
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 4804 12112 4856 12164
rect 5632 12112 5684 12164
rect 10600 12248 10652 12300
rect 12716 12248 12768 12300
rect 13912 12248 13964 12300
rect 15936 12248 15988 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 20628 12248 20680 12300
rect 21088 12248 21140 12300
rect 12532 12180 12584 12232
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 12808 12112 12860 12164
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 4988 12044 5040 12096
rect 14372 12044 14424 12096
rect 15660 12044 15712 12096
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 18972 12087 19024 12096
rect 18972 12053 18981 12087
rect 18981 12053 19015 12087
rect 19015 12053 19024 12087
rect 18972 12044 19024 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 1492 11772 1544 11824
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 8024 11704 8076 11756
rect 3148 11636 3200 11688
rect 4988 11636 5040 11688
rect 9588 11679 9640 11688
rect 3884 11611 3936 11620
rect 3884 11577 3893 11611
rect 3893 11577 3927 11611
rect 3927 11577 3936 11611
rect 3884 11568 3936 11577
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 10876 11840 10928 11892
rect 12532 11840 12584 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 10968 11679 11020 11688
rect 10968 11645 10977 11679
rect 10977 11645 11011 11679
rect 11011 11645 11020 11679
rect 10968 11636 11020 11645
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 7104 11500 7156 11552
rect 12440 11636 12492 11688
rect 14096 11772 14148 11824
rect 21640 11772 21692 11824
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 14924 11704 14976 11756
rect 15384 11704 15436 11756
rect 18236 11747 18288 11756
rect 18236 11713 18245 11747
rect 18245 11713 18279 11747
rect 18279 11713 18288 11747
rect 18236 11704 18288 11713
rect 12072 11500 12124 11552
rect 21364 11636 21416 11688
rect 21732 11636 21784 11688
rect 22008 11679 22060 11688
rect 22008 11645 22017 11679
rect 22017 11645 22051 11679
rect 22051 11645 22060 11679
rect 22008 11636 22060 11645
rect 22192 11636 22244 11688
rect 16028 11568 16080 11620
rect 16856 11568 16908 11620
rect 18604 11568 18656 11620
rect 18972 11568 19024 11620
rect 20352 11568 20404 11620
rect 15108 11500 15160 11552
rect 20628 11543 20680 11552
rect 20628 11509 20637 11543
rect 20637 11509 20671 11543
rect 20671 11509 20680 11543
rect 20628 11500 20680 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 2136 11296 2188 11348
rect 3884 11296 3936 11348
rect 4988 11228 5040 11280
rect 7564 11296 7616 11348
rect 10968 11296 11020 11348
rect 16028 11296 16080 11348
rect 20904 11296 20956 11348
rect 22100 11296 22152 11348
rect 12440 11228 12492 11280
rect 12624 11228 12676 11280
rect 15936 11271 15988 11280
rect 15936 11237 15945 11271
rect 15945 11237 15979 11271
rect 15979 11237 15988 11271
rect 15936 11228 15988 11237
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6368 11160 6420 11212
rect 7104 11160 7156 11212
rect 7472 11160 7524 11212
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 7748 11092 7800 11144
rect 14924 11160 14976 11212
rect 15752 11160 15804 11212
rect 18512 11228 18564 11280
rect 22192 11228 22244 11280
rect 10876 11092 10928 11144
rect 1860 11024 1912 11076
rect 13636 11067 13688 11076
rect 1492 10956 1544 11008
rect 13636 11033 13645 11067
rect 13645 11033 13679 11067
rect 13679 11033 13688 11067
rect 13636 11024 13688 11033
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 18420 11160 18472 11212
rect 21272 11160 21324 11212
rect 21364 11160 21416 11212
rect 22468 11203 22520 11212
rect 22468 11169 22477 11203
rect 22477 11169 22511 11203
rect 22511 11169 22520 11203
rect 22468 11160 22520 11169
rect 22652 11203 22704 11212
rect 22652 11169 22661 11203
rect 22661 11169 22695 11203
rect 22695 11169 22704 11203
rect 22652 11160 22704 11169
rect 23020 11203 23072 11212
rect 23020 11169 23029 11203
rect 23029 11169 23063 11203
rect 23063 11169 23072 11203
rect 23020 11160 23072 11169
rect 18512 11024 18564 11076
rect 21088 11024 21140 11076
rect 22008 11024 22060 11076
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 3608 10956 3660 11008
rect 3976 10956 4028 11008
rect 7012 10956 7064 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 5632 10752 5684 10804
rect 10876 10752 10928 10804
rect 3976 10616 4028 10668
rect 6920 10616 6972 10668
rect 9864 10616 9916 10668
rect 10232 10616 10284 10668
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 2044 10548 2096 10600
rect 4068 10548 4120 10600
rect 4712 10548 4764 10600
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 9680 10591 9732 10600
rect 3516 10523 3568 10532
rect 3516 10489 3525 10523
rect 3525 10489 3559 10523
rect 3559 10489 3568 10523
rect 3516 10480 3568 10489
rect 3608 10480 3660 10532
rect 2504 10412 2556 10464
rect 4620 10412 4672 10464
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 7288 10523 7340 10532
rect 7288 10489 7297 10523
rect 7297 10489 7331 10523
rect 7331 10489 7340 10523
rect 7288 10480 7340 10489
rect 7748 10480 7800 10532
rect 7472 10412 7524 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 12624 10752 12676 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14740 10795 14792 10804
rect 14740 10761 14749 10795
rect 14749 10761 14783 10795
rect 14783 10761 14792 10795
rect 14740 10752 14792 10761
rect 22100 10752 22152 10804
rect 22468 10752 22520 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 18604 10684 18656 10736
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 15384 10548 15436 10600
rect 16856 10591 16908 10600
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 19156 10591 19208 10600
rect 10324 10480 10376 10532
rect 10692 10412 10744 10464
rect 18328 10480 18380 10532
rect 19156 10557 19165 10591
rect 19165 10557 19199 10591
rect 19199 10557 19208 10591
rect 19156 10548 19208 10557
rect 20352 10591 20404 10600
rect 20352 10557 20361 10591
rect 20361 10557 20395 10591
rect 20395 10557 20404 10591
rect 20352 10548 20404 10557
rect 20536 10548 20588 10600
rect 22376 10616 22428 10668
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 17868 10412 17920 10464
rect 19432 10412 19484 10464
rect 22744 10480 22796 10532
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 3608 10208 3660 10260
rect 4804 10208 4856 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 7748 10208 7800 10260
rect 9588 10208 9640 10260
rect 5356 10183 5408 10192
rect 5356 10149 5365 10183
rect 5365 10149 5399 10183
rect 5399 10149 5408 10183
rect 5356 10140 5408 10149
rect 2044 10072 2096 10124
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3976 10072 4028 10124
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 5632 10072 5684 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6828 10115 6880 10124
rect 6368 10072 6420 10081
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 7012 10115 7064 10124
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 8208 10072 8260 10124
rect 9864 10072 9916 10124
rect 10232 10115 10284 10124
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 12348 10072 12400 10124
rect 14740 10208 14792 10260
rect 18420 10208 18472 10260
rect 18512 10208 18564 10260
rect 21364 10208 21416 10260
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 15568 10115 15620 10124
rect 12992 10004 13044 10056
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 16856 10072 16908 10124
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 22652 10115 22704 10124
rect 22652 10081 22661 10115
rect 22661 10081 22695 10115
rect 22695 10081 22704 10115
rect 22652 10072 22704 10081
rect 15016 10004 15068 10056
rect 15292 10004 15344 10056
rect 17408 10004 17460 10056
rect 2872 9936 2924 9988
rect 7656 9936 7708 9988
rect 12808 9936 12860 9988
rect 13360 9936 13412 9988
rect 17868 10004 17920 10056
rect 19156 10004 19208 10056
rect 19432 9936 19484 9988
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 7472 9868 7524 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 12900 9868 12952 9920
rect 14832 9868 14884 9920
rect 15292 9868 15344 9920
rect 15752 9911 15804 9920
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 2688 9664 2740 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 8208 9664 8260 9716
rect 15016 9664 15068 9716
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 17408 9707 17460 9716
rect 17408 9673 17417 9707
rect 17417 9673 17451 9707
rect 17451 9673 17460 9707
rect 17408 9664 17460 9673
rect 18420 9664 18472 9716
rect 20536 9664 20588 9716
rect 20628 9664 20680 9716
rect 22652 9664 22704 9716
rect 23388 9664 23440 9716
rect 18512 9596 18564 9648
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5632 9528 5684 9580
rect 7104 9528 7156 9580
rect 12256 9528 12308 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 7472 9503 7524 9512
rect 1860 9324 1912 9376
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 10140 9503 10192 9512
rect 3976 9392 4028 9444
rect 6828 9392 6880 9444
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10508 9460 10560 9512
rect 9496 9435 9548 9444
rect 9496 9401 9505 9435
rect 9505 9401 9539 9435
rect 9539 9401 9548 9435
rect 9496 9392 9548 9401
rect 10324 9392 10376 9444
rect 14924 9503 14976 9512
rect 14924 9469 14933 9503
rect 14933 9469 14967 9503
rect 14967 9469 14976 9503
rect 14924 9460 14976 9469
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 20168 9503 20220 9512
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 21272 9460 21324 9512
rect 13360 9392 13412 9444
rect 14648 9435 14700 9444
rect 14648 9401 14657 9435
rect 14657 9401 14691 9435
rect 14691 9401 14700 9435
rect 14648 9392 14700 9401
rect 15844 9435 15896 9444
rect 15844 9401 15853 9435
rect 15853 9401 15887 9435
rect 15887 9401 15896 9435
rect 15844 9392 15896 9401
rect 18236 9392 18288 9444
rect 21180 9392 21232 9444
rect 3700 9324 3752 9376
rect 5908 9324 5960 9376
rect 9680 9324 9732 9376
rect 10232 9324 10284 9376
rect 11060 9324 11112 9376
rect 15200 9324 15252 9376
rect 15568 9324 15620 9376
rect 21088 9367 21140 9376
rect 21088 9333 21097 9367
rect 21097 9333 21131 9367
rect 21131 9333 21140 9367
rect 21088 9324 21140 9333
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 21824 9324 21876 9333
rect 23112 9367 23164 9376
rect 23112 9333 23121 9367
rect 23121 9333 23155 9367
rect 23155 9333 23164 9367
rect 23112 9324 23164 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 2872 9120 2924 9172
rect 4068 9120 4120 9172
rect 5632 9120 5684 9172
rect 5908 9120 5960 9172
rect 6828 9120 6880 9172
rect 4620 9052 4672 9104
rect 9496 9120 9548 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 15016 9120 15068 9172
rect 18328 9120 18380 9172
rect 10416 9052 10468 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 5908 8984 5960 9036
rect 7656 8984 7708 9036
rect 8208 8984 8260 9036
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 17868 9052 17920 9104
rect 22284 9052 22336 9104
rect 23388 9052 23440 9104
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 14648 8984 14700 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18144 8984 18196 9036
rect 1492 8916 1544 8968
rect 3700 8916 3752 8968
rect 10324 8959 10376 8968
rect 3976 8848 4028 8900
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 12348 8916 12400 8968
rect 14096 8916 14148 8968
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 21180 8916 21232 8968
rect 21732 8959 21784 8968
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 5172 8780 5224 8832
rect 7012 8848 7064 8900
rect 11888 8848 11940 8900
rect 19248 8848 19300 8900
rect 6920 8780 6972 8832
rect 8668 8780 8720 8832
rect 10600 8780 10652 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 19432 8780 19484 8832
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 22744 8780 22796 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 1676 8576 1728 8628
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 10324 8576 10376 8628
rect 10692 8576 10744 8628
rect 12900 8576 12952 8628
rect 16672 8576 16724 8628
rect 16856 8576 16908 8628
rect 6920 8440 6972 8492
rect 7656 8440 7708 8492
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 18144 8440 18196 8492
rect 21088 8576 21140 8628
rect 21824 8440 21876 8492
rect 1860 8372 1912 8424
rect 3700 8372 3752 8424
rect 5172 8372 5224 8424
rect 6828 8372 6880 8424
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 10784 8372 10836 8424
rect 7288 8347 7340 8356
rect 7288 8313 7297 8347
rect 7297 8313 7331 8347
rect 7331 8313 7340 8347
rect 7288 8304 7340 8313
rect 7932 8304 7984 8356
rect 1676 8236 1728 8288
rect 2964 8236 3016 8288
rect 10140 8236 10192 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 11704 8236 11756 8288
rect 15844 8415 15896 8424
rect 15844 8381 15853 8415
rect 15853 8381 15887 8415
rect 15887 8381 15896 8415
rect 15844 8372 15896 8381
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 18512 8347 18564 8356
rect 18512 8313 18521 8347
rect 18521 8313 18555 8347
rect 18555 8313 18564 8347
rect 18512 8304 18564 8313
rect 19248 8304 19300 8356
rect 24492 8304 24544 8356
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 14832 8236 14884 8288
rect 16028 8279 16080 8288
rect 16028 8245 16037 8279
rect 16037 8245 16071 8279
rect 16071 8245 16080 8279
rect 16028 8236 16080 8245
rect 21732 8236 21784 8288
rect 22744 8279 22796 8288
rect 22744 8245 22753 8279
rect 22753 8245 22787 8279
rect 22787 8245 22796 8279
rect 22744 8236 22796 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 3700 8032 3752 8084
rect 3976 8032 4028 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 10784 8032 10836 8084
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 12992 8032 13044 8084
rect 19248 8032 19300 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 22376 8032 22428 8084
rect 7472 7964 7524 8016
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 4068 7896 4120 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 8760 7964 8812 8016
rect 9864 7964 9916 8016
rect 10140 8007 10192 8016
rect 10140 7973 10149 8007
rect 10149 7973 10183 8007
rect 10183 7973 10192 8007
rect 10140 7964 10192 7973
rect 10600 7964 10652 8016
rect 8208 7896 8260 7948
rect 15752 7896 15804 7948
rect 16028 7896 16080 7948
rect 16948 7896 17000 7948
rect 8668 7828 8720 7880
rect 10232 7828 10284 7880
rect 10508 7828 10560 7880
rect 18328 7896 18380 7948
rect 19432 7896 19484 7948
rect 20444 7896 20496 7948
rect 23204 7896 23256 7948
rect 18696 7828 18748 7880
rect 18972 7828 19024 7880
rect 18604 7760 18656 7812
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2228 7692 2280 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 18144 7692 18196 7744
rect 23296 7735 23348 7744
rect 23296 7701 23305 7735
rect 23305 7701 23339 7735
rect 23339 7701 23348 7735
rect 23296 7692 23348 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 23204 7531 23256 7540
rect 23204 7497 23213 7531
rect 23213 7497 23247 7531
rect 23247 7497 23256 7531
rect 23204 7488 23256 7497
rect 2228 7352 2280 7404
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 1952 7259 2004 7268
rect 1952 7225 1961 7259
rect 1961 7225 1995 7259
rect 1995 7225 2004 7259
rect 1952 7216 2004 7225
rect 3700 7148 3752 7200
rect 3792 7148 3844 7200
rect 6828 7284 6880 7336
rect 7656 7284 7708 7336
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 18512 7420 18564 7472
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 16304 7395 16356 7404
rect 9680 7284 9732 7336
rect 10140 7284 10192 7336
rect 10324 7284 10376 7336
rect 14280 7327 14332 7336
rect 7288 7216 7340 7268
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 12992 7148 13044 7200
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 16948 7352 17000 7404
rect 18604 7284 18656 7336
rect 18788 7284 18840 7336
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 17316 7216 17368 7268
rect 21732 7216 21784 7268
rect 15016 7148 15068 7200
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 2596 6944 2648 6996
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 10508 6944 10560 6996
rect 14832 6987 14884 6996
rect 14832 6953 14841 6987
rect 14841 6953 14875 6987
rect 14875 6953 14884 6987
rect 16948 6987 17000 6996
rect 14832 6944 14884 6953
rect 1952 6808 2004 6860
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 2964 6876 3016 6928
rect 5356 6876 5408 6928
rect 5816 6876 5868 6928
rect 10232 6919 10284 6928
rect 10232 6885 10241 6919
rect 10241 6885 10275 6919
rect 10275 6885 10284 6919
rect 10232 6876 10284 6885
rect 10324 6876 10376 6928
rect 11888 6919 11940 6928
rect 11888 6885 11897 6919
rect 11897 6885 11931 6919
rect 11931 6885 11940 6919
rect 11888 6876 11940 6885
rect 12348 6876 12400 6928
rect 14280 6876 14332 6928
rect 6920 6808 6972 6860
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 14004 6808 14056 6860
rect 16948 6953 16957 6987
rect 16957 6953 16991 6987
rect 16991 6953 17000 6987
rect 16948 6944 17000 6953
rect 18604 6944 18656 6996
rect 17776 6876 17828 6928
rect 16672 6808 16724 6860
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 18972 6876 19024 6928
rect 21548 6876 21600 6928
rect 18788 6851 18840 6860
rect 18788 6817 18797 6851
rect 18797 6817 18831 6851
rect 18831 6817 18840 6851
rect 18788 6808 18840 6817
rect 19892 6808 19944 6860
rect 22928 6808 22980 6860
rect 12624 6740 12676 6792
rect 15568 6740 15620 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16304 6740 16356 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 21088 6740 21140 6792
rect 21824 6783 21876 6792
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 2688 6715 2740 6724
rect 2688 6681 2697 6715
rect 2697 6681 2731 6715
rect 2731 6681 2740 6715
rect 2688 6672 2740 6681
rect 7564 6604 7616 6656
rect 19156 6647 19208 6656
rect 19156 6613 19165 6647
rect 19165 6613 19199 6647
rect 19199 6613 19208 6647
rect 19156 6604 19208 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 22008 6604 22060 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 3792 6400 3844 6452
rect 6920 6400 6972 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 17316 6443 17368 6452
rect 17316 6409 17325 6443
rect 17325 6409 17359 6443
rect 17359 6409 17368 6443
rect 17316 6400 17368 6409
rect 18144 6400 18196 6452
rect 21824 6400 21876 6452
rect 22928 6400 22980 6452
rect 23296 6400 23348 6452
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 3700 6264 3752 6316
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 3792 6196 3844 6248
rect 4988 6196 5040 6248
rect 7564 6264 7616 6316
rect 7656 6239 7708 6248
rect 5356 6128 5408 6180
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 4988 6060 5040 6112
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 8024 6239 8076 6248
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 12348 6332 12400 6384
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15568 6264 15620 6316
rect 18236 6264 18288 6316
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 20812 6264 20864 6316
rect 7932 6060 7984 6112
rect 8760 6060 8812 6112
rect 8852 6060 8904 6112
rect 9772 6196 9824 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11796 6196 11848 6248
rect 13636 6060 13688 6112
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 22836 6196 22888 6248
rect 15476 6128 15528 6180
rect 19156 6128 19208 6180
rect 20444 6171 20496 6180
rect 20444 6137 20453 6171
rect 20453 6137 20487 6171
rect 20487 6137 20496 6171
rect 20444 6128 20496 6137
rect 21088 6128 21140 6180
rect 22744 6128 22796 6180
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 2228 5856 2280 5908
rect 2412 5856 2464 5908
rect 3056 5856 3108 5908
rect 2964 5788 3016 5840
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 3608 5856 3660 5908
rect 6644 5899 6696 5908
rect 4988 5788 5040 5840
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 7656 5856 7708 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 16304 5856 16356 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 18696 5856 18748 5908
rect 19156 5856 19208 5908
rect 20812 5856 20864 5908
rect 21548 5856 21600 5908
rect 7012 5720 7064 5772
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 8024 5788 8076 5840
rect 13452 5788 13504 5840
rect 16948 5788 17000 5840
rect 18236 5788 18288 5840
rect 19892 5831 19944 5840
rect 19892 5797 19901 5831
rect 19901 5797 19935 5831
rect 19935 5797 19944 5831
rect 19892 5788 19944 5797
rect 22008 5788 22060 5840
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10416 5720 10468 5772
rect 11704 5720 11756 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 13084 5720 13136 5772
rect 14096 5720 14148 5772
rect 19064 5763 19116 5772
rect 19064 5729 19073 5763
rect 19073 5729 19107 5763
rect 19107 5729 19116 5763
rect 19064 5720 19116 5729
rect 20444 5720 20496 5772
rect 21824 5720 21876 5772
rect 22836 5763 22888 5772
rect 22836 5729 22845 5763
rect 22845 5729 22879 5763
rect 22879 5729 22888 5763
rect 22836 5720 22888 5729
rect 4620 5652 4672 5704
rect 5816 5652 5868 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7748 5584 7800 5636
rect 11244 5584 11296 5636
rect 13544 5584 13596 5636
rect 18972 5584 19024 5636
rect 21456 5584 21508 5636
rect 23572 5584 23624 5636
rect 4712 5516 4764 5568
rect 7104 5516 7156 5568
rect 8576 5516 8628 5568
rect 14096 5516 14148 5568
rect 15476 5516 15528 5568
rect 22836 5516 22888 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 4988 5312 5040 5364
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 7564 5312 7616 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 13084 5312 13136 5364
rect 21456 5355 21508 5364
rect 21456 5321 21465 5355
rect 21465 5321 21499 5355
rect 21499 5321 21508 5355
rect 21456 5312 21508 5321
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 4620 5244 4672 5296
rect 4712 5244 4764 5296
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 2044 5108 2096 5160
rect 6644 5244 6696 5296
rect 12992 5244 13044 5296
rect 6920 5176 6972 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 8760 5176 8812 5228
rect 15476 5176 15528 5228
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 8852 5108 8904 5160
rect 2596 5040 2648 5092
rect 11704 5108 11756 5160
rect 14556 5108 14608 5160
rect 19248 5176 19300 5228
rect 19524 5176 19576 5228
rect 17592 5108 17644 5160
rect 18236 5151 18288 5160
rect 18236 5117 18245 5151
rect 18245 5117 18279 5151
rect 18279 5117 18288 5151
rect 18236 5108 18288 5117
rect 21824 5151 21876 5160
rect 21824 5117 21833 5151
rect 21833 5117 21867 5151
rect 21867 5117 21876 5151
rect 21824 5108 21876 5117
rect 9956 4972 10008 5024
rect 10876 4972 10928 5024
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 14096 5040 14148 5092
rect 14188 5040 14240 5092
rect 16120 5040 16172 5092
rect 18972 5040 19024 5092
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 3608 4768 3660 4820
rect 4896 4768 4948 4820
rect 8852 4768 8904 4820
rect 12164 4768 12216 4820
rect 13636 4768 13688 4820
rect 5724 4700 5776 4752
rect 5356 4632 5408 4684
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 7472 4700 7524 4752
rect 8116 4743 8168 4752
rect 8116 4709 8125 4743
rect 8125 4709 8159 4743
rect 8159 4709 8168 4743
rect 8116 4700 8168 4709
rect 13544 4743 13596 4752
rect 13544 4709 13553 4743
rect 13553 4709 13587 4743
rect 13587 4709 13596 4743
rect 13544 4700 13596 4709
rect 6000 4632 6052 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 8576 4675 8628 4684
rect 6460 4632 6512 4641
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 11152 4632 11204 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 7472 4564 7524 4616
rect 18972 4768 19024 4820
rect 20812 4768 20864 4820
rect 21824 4768 21876 4820
rect 19616 4700 19668 4752
rect 19984 4700 20036 4752
rect 22836 4743 22888 4752
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 16856 4632 16908 4684
rect 17592 4632 17644 4684
rect 19064 4675 19116 4684
rect 19064 4641 19073 4675
rect 19073 4641 19107 4675
rect 19107 4641 19116 4675
rect 19064 4632 19116 4641
rect 19432 4632 19484 4684
rect 22468 4632 22520 4684
rect 23572 4632 23624 4684
rect 15752 4607 15804 4616
rect 8484 4496 8536 4548
rect 12624 4496 12676 4548
rect 14280 4496 14332 4548
rect 3700 4428 3752 4480
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 5356 4428 5408 4437
rect 6920 4428 6972 4480
rect 13360 4428 13412 4480
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 16304 4564 16356 4616
rect 21640 4564 21692 4616
rect 16948 4428 17000 4480
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 19984 4428 20036 4480
rect 20628 4428 20680 4480
rect 21916 4428 21968 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 2596 4267 2648 4276
rect 2596 4233 2605 4267
rect 2605 4233 2639 4267
rect 2639 4233 2648 4267
rect 2596 4224 2648 4233
rect 5540 4224 5592 4276
rect 6460 4224 6512 4276
rect 4804 4156 4856 4208
rect 5356 4156 5408 4208
rect 7104 4156 7156 4208
rect 7288 4224 7340 4276
rect 9864 4224 9916 4276
rect 10876 4267 10928 4276
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 16856 4224 16908 4276
rect 17592 4267 17644 4276
rect 17592 4233 17601 4267
rect 17601 4233 17635 4267
rect 17635 4233 17644 4267
rect 17592 4224 17644 4233
rect 22468 4267 22520 4276
rect 22468 4233 22477 4267
rect 22477 4233 22511 4267
rect 22511 4233 22520 4267
rect 22468 4224 22520 4233
rect 23572 4224 23624 4276
rect 15752 4156 15804 4208
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 12164 4088 12216 4140
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 13452 4088 13504 4140
rect 13912 4088 13964 4140
rect 14556 4088 14608 4140
rect 14740 4088 14792 4140
rect 3148 3952 3200 4004
rect 3700 3952 3752 4004
rect 5448 3952 5500 4004
rect 9220 3995 9272 4004
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 9220 3961 9229 3995
rect 9229 3961 9263 3995
rect 9263 3961 9272 3995
rect 9220 3952 9272 3961
rect 8484 3884 8536 3936
rect 9588 3884 9640 3936
rect 14280 4020 14332 4072
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 19984 4088 20036 4140
rect 21916 4131 21968 4140
rect 15844 4020 15896 4072
rect 16120 4063 16172 4072
rect 16120 4029 16129 4063
rect 16129 4029 16163 4063
rect 16163 4029 16172 4063
rect 16120 4020 16172 4029
rect 11336 3884 11388 3936
rect 13360 3952 13412 4004
rect 14188 3952 14240 4004
rect 14924 3952 14976 4004
rect 17960 4020 18012 4072
rect 19616 4063 19668 4072
rect 17408 3884 17460 3936
rect 19616 4029 19625 4063
rect 19625 4029 19659 4063
rect 19659 4029 19668 4063
rect 19616 4020 19668 4029
rect 20352 4020 20404 4072
rect 21456 4063 21508 4072
rect 21456 4029 21465 4063
rect 21465 4029 21499 4063
rect 21499 4029 21508 4063
rect 21456 4020 21508 4029
rect 21640 4063 21692 4072
rect 21640 4029 21649 4063
rect 21649 4029 21683 4063
rect 21683 4029 21692 4063
rect 21640 4020 21692 4029
rect 21916 4097 21925 4131
rect 21925 4097 21959 4131
rect 21959 4097 21968 4131
rect 21916 4088 21968 4097
rect 22008 4063 22060 4072
rect 22008 4029 22017 4063
rect 22017 4029 22051 4063
rect 22051 4029 22060 4063
rect 22008 4020 22060 4029
rect 19248 3952 19300 4004
rect 20904 3952 20956 4004
rect 20444 3884 20496 3936
rect 22652 3884 22704 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 3700 3680 3752 3732
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 12900 3680 12952 3732
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 5448 3612 5500 3664
rect 10600 3612 10652 3664
rect 11520 3612 11572 3664
rect 14556 3612 14608 3664
rect 5264 3544 5316 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 6000 3544 6052 3596
rect 7104 3544 7156 3596
rect 11888 3544 11940 3596
rect 13912 3544 13964 3596
rect 14188 3587 14240 3596
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 16120 3612 16172 3664
rect 17684 3612 17736 3664
rect 21824 3612 21876 3664
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 13728 3476 13780 3528
rect 16304 3544 16356 3596
rect 16948 3587 17000 3596
rect 16948 3553 16957 3587
rect 16957 3553 16991 3587
rect 16991 3553 17000 3587
rect 16948 3544 17000 3553
rect 19064 3544 19116 3596
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 20904 3476 20956 3528
rect 21088 3519 21140 3528
rect 21088 3485 21097 3519
rect 21097 3485 21131 3519
rect 21131 3485 21140 3519
rect 21088 3476 21140 3485
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21456 3476 21508 3528
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 8576 3340 8628 3392
rect 8852 3383 8904 3392
rect 8852 3349 8861 3383
rect 8861 3349 8895 3383
rect 8895 3349 8904 3383
rect 8852 3340 8904 3349
rect 14740 3340 14792 3392
rect 19984 3340 20036 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 8852 3136 8904 3188
rect 11520 3136 11572 3188
rect 12900 3179 12952 3188
rect 12900 3145 12909 3179
rect 12909 3145 12943 3179
rect 12943 3145 12952 3179
rect 12900 3136 12952 3145
rect 13636 3136 13688 3188
rect 16304 3136 16356 3188
rect 16948 3136 17000 3188
rect 17684 3136 17736 3188
rect 20352 3136 20404 3188
rect 8116 3111 8168 3120
rect 1584 3000 1636 3052
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 5724 3000 5776 3052
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 10232 3068 10284 3120
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 2596 2907 2648 2916
rect 296 2796 348 2848
rect 2596 2873 2605 2907
rect 2605 2873 2639 2907
rect 2639 2873 2648 2907
rect 2596 2864 2648 2873
rect 2688 2796 2740 2848
rect 5448 2975 5500 2984
rect 5172 2907 5224 2916
rect 5172 2873 5181 2907
rect 5181 2873 5215 2907
rect 5215 2873 5224 2907
rect 5172 2864 5224 2873
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 7564 2932 7616 2984
rect 9220 2932 9272 2984
rect 11244 2975 11296 2984
rect 9772 2864 9824 2916
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 11980 2975 12032 2984
rect 11980 2941 11989 2975
rect 11989 2941 12023 2975
rect 12023 2941 12032 2975
rect 11980 2932 12032 2941
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 17224 3000 17276 3052
rect 19432 3043 19484 3052
rect 19432 3009 19441 3043
rect 19441 3009 19475 3043
rect 19475 3009 19484 3043
rect 19432 3000 19484 3009
rect 21364 3111 21416 3120
rect 21364 3077 21373 3111
rect 21373 3077 21407 3111
rect 21407 3077 21416 3111
rect 21364 3068 21416 3077
rect 21824 3136 21876 3188
rect 22652 3179 22704 3188
rect 22652 3145 22661 3179
rect 22661 3145 22695 3179
rect 22695 3145 22704 3179
rect 22652 3136 22704 3145
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 15476 2932 15528 2984
rect 12072 2864 12124 2916
rect 4712 2796 4764 2848
rect 6000 2796 6052 2848
rect 10140 2796 10192 2848
rect 11336 2796 11388 2848
rect 14372 2796 14424 2848
rect 15292 2796 15344 2848
rect 20444 2975 20496 2984
rect 20444 2941 20453 2975
rect 20453 2941 20487 2975
rect 20487 2941 20496 2975
rect 20444 2932 20496 2941
rect 20628 2932 20680 2984
rect 22008 2932 22060 2984
rect 19892 2864 19944 2916
rect 21088 2864 21140 2916
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 2596 2592 2648 2644
rect 4712 2592 4764 2644
rect 5172 2592 5224 2644
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12624 2592 12676 2644
rect 13728 2635 13780 2644
rect 4988 2524 5040 2576
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 14188 2592 14240 2644
rect 14372 2524 14424 2576
rect 12900 2456 12952 2508
rect 15476 2592 15528 2644
rect 17684 2592 17736 2644
rect 19064 2635 19116 2644
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 21364 2635 21416 2644
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 21456 2592 21508 2644
rect 14740 2567 14792 2576
rect 14740 2533 14749 2567
rect 14749 2533 14783 2567
rect 14783 2533 14792 2567
rect 14740 2524 14792 2533
rect 18972 2388 19024 2440
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 12164 1300 12216 1352
rect 22376 1300 22428 1352
rect 4896 8 4948 60
rect 15200 8 15252 60
<< metal2 >>
rect 938 27282 994 27971
rect 3422 27282 3478 27971
rect 5906 27282 5962 27971
rect 938 27254 1164 27282
rect 938 27171 994 27254
rect 1136 12306 1164 27254
rect 3344 27254 3478 27282
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1674 25120 1730 25129
rect 1674 25055 1730 25064
rect 1688 24274 1716 25055
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1688 23866 1716 24210
rect 2056 24206 2084 25230
rect 3344 24342 3372 27254
rect 3422 27171 3478 27254
rect 5552 27254 5962 27282
rect 5552 25362 5580 27254
rect 5906 27171 5962 27254
rect 8390 27260 8446 27971
rect 10874 27282 10930 27971
rect 13358 27282 13414 27971
rect 8390 27208 8392 27260
rect 8444 27208 8446 27260
rect 8390 27171 8446 27208
rect 10612 27254 10930 27282
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 5540 25356 5592 25362
rect 5540 25298 5592 25304
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 5000 24954 5028 25298
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 5184 24750 5212 25094
rect 7300 24954 7328 25230
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 8300 24948 8352 24954
rect 8300 24890 8352 24896
rect 7300 24750 7328 24890
rect 5172 24744 5224 24750
rect 5172 24686 5224 24692
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 5356 24608 5408 24614
rect 5356 24550 5408 24556
rect 3332 24336 3384 24342
rect 3332 24278 3384 24284
rect 4724 24274 4752 24550
rect 5368 24274 5396 24550
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1872 23186 1900 24006
rect 2056 23866 2084 24142
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 2976 23662 3004 24142
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3160 23662 3188 24006
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2964 23656 3016 23662
rect 2964 23598 3016 23604
rect 3148 23656 3200 23662
rect 3148 23598 3200 23604
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1860 23180 1912 23186
rect 1860 23122 1912 23128
rect 1596 22234 1624 23122
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 2136 22976 2188 22982
rect 2136 22918 2188 22924
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 1214 21448 1270 21457
rect 1214 21383 1270 21392
rect 1124 12300 1176 12306
rect 1124 12242 1176 12248
rect 1228 9625 1256 21383
rect 1688 21078 1716 22918
rect 2148 22574 2176 22918
rect 2424 22642 2452 23530
rect 2608 23322 2636 23598
rect 4632 23594 4660 24210
rect 4724 23798 4752 24210
rect 4988 24132 5040 24138
rect 4988 24074 5040 24080
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 4620 23588 4672 23594
rect 4620 23530 4672 23536
rect 4632 23474 4660 23530
rect 4448 23446 4660 23474
rect 4448 23322 4476 23446
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 5000 23254 5028 24074
rect 5184 23730 5212 24210
rect 5368 23866 5396 24210
rect 6380 23866 6408 24686
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 6368 23860 6420 23866
rect 6368 23802 6420 23808
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5920 23322 5948 23802
rect 6380 23662 6408 23802
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 6380 23254 6408 23598
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5724 23248 5776 23254
rect 5724 23190 5776 23196
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2884 22506 2912 23054
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2596 22092 2648 22098
rect 2596 22034 2648 22040
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1676 21072 1728 21078
rect 1676 21014 1728 21020
rect 1688 20942 1716 21014
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1688 19310 1716 20878
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 2056 20398 2084 20742
rect 2148 20602 2176 21422
rect 2332 21418 2360 21966
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2516 21554 2544 21830
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2240 21010 2268 21286
rect 2332 21010 2360 21354
rect 2516 21010 2544 21490
rect 2608 21486 2636 22034
rect 2884 21690 2912 22442
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 3620 21146 3648 22918
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 5000 22778 5028 23190
rect 5736 22778 5764 23190
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4172 22234 4200 22442
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4160 22228 4212 22234
rect 4160 22170 4212 22176
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4632 21350 4660 22374
rect 5724 22160 5776 22166
rect 5724 22102 5776 22108
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5368 21690 5396 22034
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2504 21004 2556 21010
rect 2504 20946 2556 20952
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1688 18834 1716 19246
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 2056 18290 2084 20334
rect 2148 19922 2176 20538
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 18902 2176 19858
rect 2240 19310 2268 20946
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2332 18970 2360 20946
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 2424 20466 2452 20810
rect 2412 20460 2464 20466
rect 2412 20402 2464 20408
rect 2412 19984 2464 19990
rect 2516 19972 2544 20946
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3528 20398 3556 20810
rect 3620 20806 3648 21082
rect 4632 21010 4660 21286
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3528 20058 3556 20334
rect 4632 20262 4660 20946
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 2464 19944 2544 19972
rect 2412 19926 2464 19932
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 19514 3556 19654
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3528 19310 3556 19450
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 4080 19242 4108 19858
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2056 17814 2084 18226
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 16726 1716 17478
rect 2056 17134 2084 17750
rect 2424 17202 2452 19110
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16046 1716 16390
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15502 1716 15982
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15366 1716 15438
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 14074 1716 15302
rect 1872 14618 1900 15506
rect 2056 14958 2084 17070
rect 2320 16720 2372 16726
rect 2320 16662 2372 16668
rect 2332 16046 2360 16662
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2228 15564 2280 15570
rect 2332 15552 2360 15982
rect 2516 15570 2544 16526
rect 2608 15978 2636 18090
rect 2976 17882 3004 18090
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3068 17814 3096 18770
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 3160 17066 3188 18566
rect 4080 18290 4108 19178
rect 4632 18698 4660 20198
rect 4816 19922 4844 20198
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 5368 19514 5396 21626
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5368 18902 5396 19450
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4816 18358 4844 18566
rect 5092 18426 5120 18770
rect 5644 18766 5672 21558
rect 5736 21078 5764 22102
rect 6104 22098 6132 22918
rect 7208 22778 7236 23122
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6104 21622 6132 22034
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 5724 21072 5776 21078
rect 6092 21072 6144 21078
rect 5724 21014 5776 21020
rect 5828 21032 6092 21060
rect 5736 20602 5764 21014
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5828 20262 5856 21032
rect 6092 21014 6144 21020
rect 6092 20936 6144 20942
rect 6196 20924 6224 22374
rect 6144 20896 6224 20924
rect 6092 20878 6144 20884
rect 6104 20398 6132 20878
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5736 19310 5764 19790
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18970 5764 19246
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 5368 18290 5396 18702
rect 5736 18426 5764 18906
rect 5828 18426 5856 20198
rect 6104 19922 6132 20334
rect 6828 19984 6880 19990
rect 6828 19926 6880 19932
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6380 19514 6408 19790
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6288 18834 6316 19246
rect 6380 18970 6408 19450
rect 6840 18970 6868 19926
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 7116 18902 7144 19246
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 6288 18358 6316 18770
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16794 3188 17002
rect 3252 16794 3280 17682
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3712 16794 3740 17002
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 4080 16454 4108 17070
rect 4632 16998 4660 17682
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 5000 16658 5028 17478
rect 5368 17134 5396 17614
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16114 4108 16390
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 4908 15638 4936 16458
rect 5000 16250 5028 16594
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 2504 15564 2556 15570
rect 2280 15524 2360 15552
rect 2424 15524 2504 15552
rect 2228 15506 2280 15512
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 2424 14906 2452 15524
rect 2504 15506 2556 15512
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2516 15026 2544 15370
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2056 13938 2084 14894
rect 2424 14878 2544 14906
rect 2516 14414 2544 14878
rect 2608 14482 2636 15574
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4908 15162 4936 15574
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 3620 14958 3648 15030
rect 5092 14958 5120 16934
rect 5368 16046 5396 17070
rect 5460 16658 5488 17274
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 6104 16658 6132 17002
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5460 15366 5488 16594
rect 5920 16114 5948 16594
rect 6104 16250 6132 16594
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6104 16046 6132 16186
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6656 15978 6684 17070
rect 6840 16794 6868 17682
rect 6932 17338 6960 17682
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7484 16114 7512 17614
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6656 15638 6684 15914
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 3620 14618 3648 14894
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 4356 14482 4384 14826
rect 5552 14822 5580 15574
rect 7208 15502 7236 15982
rect 7484 15706 7512 16050
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6288 15162 6316 15438
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13190 2176 13806
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1596 12764 1624 13126
rect 2148 12850 2176 13126
rect 2424 12986 2452 14350
rect 2608 13530 2636 14418
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 1676 12776 1728 12782
rect 1596 12736 1676 12764
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 11830 1532 12174
rect 1492 11824 1544 11830
rect 1492 11766 1544 11772
rect 1504 11014 1532 11766
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1214 9616 1270 9625
rect 1214 9551 1270 9560
rect 1504 8974 1532 10950
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 7732 1532 8910
rect 1596 7857 1624 12736
rect 1676 12718 1728 12724
rect 2608 12442 2636 13466
rect 2700 12986 2728 13874
rect 2792 13394 2820 14282
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 5000 14074 5028 14418
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2976 13530 3004 13738
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 4080 13462 4108 13806
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2792 12646 2820 13330
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3620 12714 3648 13126
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4632 12986 4660 13330
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12918 4752 13738
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 13258 5212 13330
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12986 5212 13194
rect 5552 12986 5580 14758
rect 5644 14618 5672 14894
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5644 13870 5672 14554
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6288 13938 6316 14214
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12442 2820 12582
rect 5368 12442 5396 12718
rect 6932 12714 6960 13874
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 1688 11898 1716 12242
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 2148 11354 2176 12174
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3160 11694 3188 12038
rect 3620 11762 3648 12038
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10606 1900 11018
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 1674 10432 1730 10441
rect 1674 10367 1730 10376
rect 1688 9042 1716 10367
rect 2056 10130 2084 10542
rect 2516 10470 2544 11494
rect 3620 11098 3648 11698
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 11354 3924 11562
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3620 11070 3740 11098
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10130 2544 10406
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 9722 2728 10066
rect 2884 9994 2912 10950
rect 3620 10538 3648 10950
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1688 8634 1716 8978
rect 1872 8838 1900 9318
rect 2884 9178 2912 9930
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9586 3004 9862
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1872 8430 1900 8774
rect 3528 8634 3556 10474
rect 3620 10266 3648 10474
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3712 9382 3740 11070
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10674 4016 10950
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 10130 4016 10610
rect 4816 10606 4844 12106
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11694 5028 12038
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 11286 5028 11630
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 8974 3740 9318
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3712 8430 3740 8910
rect 3988 8906 4016 9386
rect 4080 9178 4108 10542
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4632 9110 4660 10406
rect 4724 10130 4752 10542
rect 4816 10266 4844 10542
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9586 4752 10066
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 5092 9042 5120 12242
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11762 5672 12106
rect 7024 11898 7052 15438
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13394 7236 14214
rect 7484 14074 7512 14418
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13530 7328 13738
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7116 12986 7144 13330
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7392 12782 7420 13874
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7484 12918 7512 13330
rect 7576 13190 7604 24686
rect 8036 24410 8064 24686
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7668 23662 7696 24210
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 7760 23662 7788 24142
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7748 23656 7800 23662
rect 7748 23598 7800 23604
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 7668 21078 7696 23598
rect 8128 23322 8156 23598
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8312 23186 8340 24890
rect 8404 24614 8432 25298
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 8496 23866 8524 24210
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 8588 23186 8616 25094
rect 9416 24818 9444 25094
rect 10428 24818 10456 25094
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 8772 23662 8800 24142
rect 9416 24138 9444 24754
rect 10612 24750 10640 27254
rect 10874 27171 10930 27254
rect 11704 27260 11756 27266
rect 11704 27202 11756 27208
rect 13096 27254 13414 27282
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10888 24750 10916 25094
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9416 23866 9444 24074
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 9876 23186 9904 24618
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7944 22234 7972 22374
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7852 20398 7880 21082
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 19514 7880 20334
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 8128 19310 8156 19790
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7852 18222 7880 18770
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 8036 16794 8064 18022
rect 8220 17746 8248 22918
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8404 22098 8432 22510
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8404 21690 8432 22034
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8496 20466 8524 22442
rect 8588 22234 8616 23122
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 9968 22438 9996 22918
rect 10520 22710 10548 22918
rect 10888 22778 10916 24686
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10980 23798 11008 24210
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10508 22704 10560 22710
rect 10508 22646 10560 22652
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10232 22500 10284 22506
rect 10232 22442 10284 22448
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8588 21146 8616 21422
rect 8864 21146 8892 22374
rect 9968 22030 9996 22374
rect 10244 22098 10272 22442
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9692 21554 9720 21898
rect 10428 21554 10456 22578
rect 10520 22098 10548 22646
rect 10980 22574 11008 22918
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8588 20330 8616 20810
rect 10152 20602 10180 21354
rect 10428 21010 10456 21490
rect 10520 21078 10548 22034
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10428 20534 10456 20946
rect 10416 20528 10468 20534
rect 10416 20470 10468 20476
rect 8576 20324 8628 20330
rect 8576 20266 8628 20272
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 8588 19514 8616 20266
rect 9876 19922 9904 20266
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9324 19718 9352 19858
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 9324 18970 9352 19654
rect 9876 19378 9904 19858
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 10336 19242 10364 19654
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17882 8340 18022
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 16998 8616 17682
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 15978 8064 16730
rect 8588 16658 8616 16934
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8496 15026 8524 16050
rect 8588 15706 8616 16594
rect 8772 16454 8800 18226
rect 10060 18222 10088 19110
rect 10336 18630 10364 19178
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18426 10364 18566
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9048 16998 9076 17682
rect 9876 17542 9904 18158
rect 10060 17882 10088 18158
rect 10336 18154 10364 18362
rect 10520 18222 10548 18906
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9324 17134 9352 17478
rect 10060 17134 10088 17818
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7668 13462 7696 14758
rect 7852 14464 7880 14826
rect 8496 14618 8524 14962
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 7932 14476 7984 14482
rect 7852 14436 7932 14464
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 13938 7788 14350
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7748 13388 7800 13394
rect 7852 13376 7880 14436
rect 7932 14418 7984 14424
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 13462 7972 13738
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 8036 13394 8064 14282
rect 7800 13348 7880 13376
rect 8024 13388 8076 13394
rect 7748 13330 7800 13336
rect 8024 13330 8076 13336
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 12442 7420 12718
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7012 11892 7064 11898
rect 6932 11852 7012 11880
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 5644 10810 5672 11154
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5368 9722 5396 10134
rect 5644 10130 5672 10746
rect 6380 10130 6408 11154
rect 6932 10674 6960 11852
rect 7012 11834 7064 11840
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11218 7144 11494
rect 7576 11354 7604 13126
rect 7760 12442 7788 13330
rect 8036 12850 8064 13330
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8220 12442 8248 12922
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11762 8064 12242
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5644 9586 5672 10066
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5644 9178 5672 9522
rect 6840 9450 6868 10066
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 6840 9178 6868 9386
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 1676 8288 1728 8294
rect 1676 8230 1728 8236
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 1582 7848 1638 7857
rect 1582 7783 1638 7792
rect 1584 7744 1636 7750
rect 1504 7704 1584 7732
rect 1584 7686 1636 7692
rect 1596 3058 1624 7686
rect 1688 6798 1716 8230
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 7410 2268 7686
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1964 6866 1992 7210
rect 2240 6866 2268 7346
rect 2424 7342 2452 7890
rect 2976 7342 3004 8230
rect 3712 8090 3740 8366
rect 3988 8090 4016 8842
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 5092 8090 5120 8978
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8430 5212 8774
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5920 8090 5948 8978
rect 6932 8838 6960 10610
rect 7024 10130 7052 10950
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 10266 7328 10474
rect 7484 10470 7512 11154
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7760 10538 7788 11086
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 9568 7052 10066
rect 7484 9926 7512 10406
rect 7760 10266 7788 10474
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7104 9580 7156 9586
rect 7024 9540 7104 9568
rect 7024 8906 7052 9540
rect 7104 9522 7156 9528
rect 7484 9518 7512 9862
rect 7668 9518 7696 9930
rect 8220 9722 8248 10066
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 9042 7696 9454
rect 8220 9042 8248 9658
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8498 6960 8774
rect 7668 8498 7696 8978
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6840 7954 6868 8366
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 4080 7342 4108 7890
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 2608 7002 2636 7278
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1688 5166 1716 6734
rect 1676 5160 1728 5166
rect 1964 5148 1992 6802
rect 2240 5914 2268 6802
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5914 2452 6190
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2608 5778 2636 6938
rect 2976 6934 3004 7278
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2700 6322 2728 6666
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2976 5846 3004 6870
rect 3620 5914 3648 6938
rect 3712 6322 3740 7142
rect 3804 6458 3832 7142
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3804 6254 3832 6394
rect 5000 6254 5028 7142
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 3792 6248 3844 6254
rect 4988 6248 5040 6254
rect 3792 6190 3844 6196
rect 4908 6208 4988 6236
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2044 5160 2096 5166
rect 1964 5120 2044 5148
rect 1676 5102 1728 5108
rect 2044 5102 2096 5108
rect 1688 4826 1716 5102
rect 2056 4826 2084 5102
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2608 4282 2636 5034
rect 3068 4826 3096 5850
rect 3620 4826 3648 5850
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4632 5302 4660 5646
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5302 4752 5510
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4908 4826 4936 6208
rect 4988 6190 5040 6196
rect 5368 6186 5396 6870
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5000 5846 5028 6054
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5000 5370 5028 5782
rect 5368 5370 5396 6122
rect 5828 5710 5856 6870
rect 6656 5914 6684 7686
rect 6840 7342 6868 7890
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 7300 7274 7328 8298
rect 7944 8090 7972 8298
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 7546 7512 7958
rect 8220 7954 8248 8978
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 6458 6960 6802
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 6656 5302 6684 5850
rect 6932 5710 6960 6394
rect 7576 6322 7604 6598
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 5778 7052 6122
rect 7576 5778 7604 6258
rect 7668 6254 7696 7278
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5914 7696 6190
rect 7944 6118 7972 6802
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 8036 5846 8064 6190
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6932 5234 6960 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 3068 4154 3096 4762
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 4486 5396 4626
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 3068 4126 3188 4154
rect 3160 4010 3188 4126
rect 3712 4010 3740 4422
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 5368 4214 5396 4422
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3712 3738 3740 3946
rect 4816 3738 4844 4150
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 5460 3670 5488 3946
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5264 3596 5316 3602
rect 5184 3556 5264 3584
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 296 2848 348 2854
rect 296 2790 348 2796
rect 18 82 74 800
rect 308 82 336 2790
rect 2056 2650 2084 2994
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2608 2650 2636 2858
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 18 54 336 82
rect 2410 82 2466 800
rect 2700 82 2728 2790
rect 4724 2650 4752 2790
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5000 2582 5028 3470
rect 5184 2922 5212 3556
rect 5264 3538 5316 3544
rect 5460 2990 5488 3606
rect 5552 3602 5580 4218
rect 5736 3942 5764 4694
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3602 5764 3878
rect 6012 3602 6040 4626
rect 6472 4282 6500 4626
rect 6932 4486 6960 5170
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7116 4298 7144 5510
rect 7576 5370 7604 5714
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7760 5234 7788 5578
rect 8588 5574 8616 14894
rect 8772 14822 8800 16390
rect 9048 15026 9076 16934
rect 9324 16794 9352 17070
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9876 16250 9904 16594
rect 10244 16454 10272 16934
rect 10796 16726 10824 17002
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 9864 16244 9916 16250
rect 9784 16204 9864 16232
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9692 13938 9720 14418
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9220 13864 9272 13870
rect 9784 13814 9812 16204
rect 9864 16186 9916 16192
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14482 10088 14758
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9220 13806 9272 13812
rect 9232 13530 9260 13806
rect 9692 13786 9812 13814
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9600 10266 9628 11630
rect 9692 10606 9720 13786
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9784 12646 9812 13398
rect 9876 13326 9904 14282
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9876 12714 9904 13262
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12442 9812 12582
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 10674 9904 11154
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9876 10130 9904 10406
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9178 9536 9386
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 7886 8708 8774
rect 9692 8430 9720 9318
rect 9968 9178 9996 9862
rect 10152 9518 10180 15982
rect 10244 15570 10272 16390
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10244 15162 10272 15506
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10428 15065 10456 15914
rect 10796 15706 10824 16662
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10414 15056 10470 15065
rect 10414 14991 10470 15000
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10244 14074 10272 14214
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10612 13462 10640 15302
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10704 14006 10732 14418
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10612 12986 10640 13398
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12306 10640 12582
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10888 11898 10916 22374
rect 10980 22098 11008 22510
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 11072 18714 11100 24754
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11440 23866 11468 24210
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11532 23322 11560 24618
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11256 22574 11284 22986
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11256 22166 11284 22510
rect 11624 22234 11652 23802
rect 11612 22228 11664 22234
rect 11612 22170 11664 22176
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11440 20262 11468 20946
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11164 19310 11192 19790
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11164 18970 11192 19246
rect 11440 19174 11468 20198
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 19378 11560 19858
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11532 19242 11560 19314
rect 11520 19236 11572 19242
rect 11520 19178 11572 19184
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 10980 18358 11008 18702
rect 11072 18686 11192 18714
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10968 18352 11020 18358
rect 10968 18294 11020 18300
rect 11072 17542 11100 18566
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11072 16590 11100 17478
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 15910 11100 16526
rect 11164 16114 11192 18686
rect 11440 18630 11468 19110
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11440 17746 11468 18566
rect 11716 17746 11744 27202
rect 12624 25356 12676 25362
rect 12624 25298 12676 25304
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 21690 12020 24006
rect 12268 23798 12296 24210
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12268 23322 12296 23734
rect 12360 23594 12388 24006
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 12360 21146 12388 23530
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22778 12480 23054
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12544 22012 12572 23598
rect 12636 23186 12664 25298
rect 13096 24614 13124 27254
rect 13358 27171 13414 27254
rect 15842 27282 15898 27971
rect 18326 27282 18382 27971
rect 20810 27282 20866 27971
rect 23294 27282 23350 27971
rect 25686 27282 25742 27971
rect 15842 27254 15976 27282
rect 15842 27171 15898 27254
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13188 24818 13216 25298
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 13556 24274 13584 25094
rect 14200 24750 14228 25162
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14476 24750 14504 25094
rect 15948 24750 15976 27254
rect 18064 27254 18382 27282
rect 16120 25356 16172 25362
rect 16120 25298 16172 25304
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16132 24954 16160 25298
rect 16776 24954 16804 25298
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16120 24948 16172 24954
rect 16764 24948 16816 24954
rect 16120 24890 16172 24896
rect 16684 24908 16764 24936
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 14200 24410 14228 24686
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14476 24342 14504 24686
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12820 23322 12848 24142
rect 12900 24132 12952 24138
rect 12900 24074 12952 24080
rect 12912 23730 12940 24074
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12636 22166 12664 23122
rect 13464 23118 13492 24210
rect 13556 23866 13584 24210
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13556 23186 13584 23802
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 14660 23050 14688 23530
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 12624 22024 12676 22030
rect 12544 21984 12624 22012
rect 12624 21966 12676 21972
rect 12636 21486 12664 21966
rect 13004 21554 13032 22034
rect 13188 22030 13216 22646
rect 14936 22642 14964 24618
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15488 23730 15516 24346
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15672 23662 15700 24278
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16132 23662 16160 23734
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15028 22642 15056 22918
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 14016 22234 14044 22442
rect 15304 22234 15332 22442
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 13004 21078 13032 21490
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13372 21146 13400 21354
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 14200 21010 14228 22034
rect 15948 22030 15976 23054
rect 16040 22642 16068 23530
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16224 23118 16252 23462
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16224 22778 16252 23054
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16316 22574 16344 24210
rect 16684 24206 16712 24908
rect 16764 24890 16816 24896
rect 16960 24274 16988 25094
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17328 24410 17356 24550
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16684 23866 16712 24142
rect 16776 23866 16804 24210
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16396 23792 16448 23798
rect 16396 23734 16448 23740
rect 16408 23322 16436 23734
rect 16684 23474 16712 23802
rect 16776 23662 16804 23802
rect 16960 23798 16988 24210
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16592 23446 16712 23474
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16592 23118 16620 23446
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 14752 21146 14780 21966
rect 16316 21690 16344 22510
rect 16776 22234 16804 23190
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 17880 22098 17908 22510
rect 18064 22506 18092 27254
rect 18326 27171 18382 27254
rect 20732 27254 20866 27282
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18524 23322 18552 24074
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18524 22778 18552 23258
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14740 21140 14792 21146
rect 14660 21100 14740 21128
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13740 20262 13768 20334
rect 13832 20262 13860 20946
rect 14660 20466 14688 21100
rect 14740 21082 14792 21088
rect 14936 21010 14964 21286
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14004 20460 14056 20466
rect 14648 20460 14700 20466
rect 14056 20420 14136 20448
rect 14004 20402 14056 20408
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13004 19922 13032 20198
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 18834 12112 19654
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18902 12756 19178
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 17882 12112 18770
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11440 16998 11468 17682
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11532 16726 11560 17478
rect 12084 16998 12112 17614
rect 12912 17202 12940 19246
rect 13004 18630 13032 19858
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14016 18630 14044 19246
rect 14108 18970 14136 20420
rect 14648 20402 14700 20408
rect 14752 20330 14780 20810
rect 16316 20466 16344 21626
rect 16592 21350 16620 22034
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18156 21690 18184 21966
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16960 21010 16988 21354
rect 18156 21078 18184 21626
rect 18616 21622 18644 22102
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18340 21146 18368 21422
rect 18604 21412 18656 21418
rect 18604 21354 18656 21360
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16500 20602 16528 20946
rect 16960 20602 16988 20946
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 16488 20596 16540 20602
rect 16488 20538 16540 20544
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 14280 20324 14332 20330
rect 14280 20266 14332 20272
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 14292 19242 14320 20266
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19718 14504 20198
rect 14752 20058 14780 20266
rect 16500 20058 16528 20538
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16960 19990 16988 20538
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 17788 19922 17816 20878
rect 18340 19922 18368 21082
rect 18616 20806 18644 21354
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 19310 14504 19654
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17814 13124 18022
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13280 17338 13308 17682
rect 14016 17678 14044 18566
rect 14108 18290 14136 18906
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11532 16250 11560 16662
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 14414 11100 15846
rect 11164 15706 11192 16050
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 12084 15201 12112 16934
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14006 11376 14350
rect 11808 14074 11836 14486
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13462 11928 13874
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 12544 12238 12572 15642
rect 12820 14958 12848 16526
rect 12912 16250 12940 17138
rect 14016 17134 14044 17614
rect 14476 17270 14504 19246
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14752 17270 14780 18090
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14936 17134 14964 17750
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 13188 16454 13216 17070
rect 14016 16794 14044 17070
rect 14108 16794 14136 17070
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14844 16794 14872 17002
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15120 16658 15148 18226
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 13188 16046 13216 16390
rect 15120 16250 15148 16594
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13096 15026 13124 15506
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 15026 13584 15302
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 13870 12756 14758
rect 13096 14600 13124 14962
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13176 14612 13228 14618
rect 13096 14572 13176 14600
rect 13176 14554 13228 14560
rect 13372 13870 13400 14894
rect 13556 13870 13584 14962
rect 14200 14482 14228 15846
rect 14832 15428 14884 15434
rect 14832 15370 14884 15376
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 14958 14596 15302
rect 14844 15201 14872 15370
rect 14830 15192 14886 15201
rect 14830 15127 14886 15136
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 12716 13864 12768 13870
rect 12900 13864 12952 13870
rect 12716 13806 12768 13812
rect 12820 13824 12900 13852
rect 12728 13462 12756 13806
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12442 12664 12650
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11898 12572 12174
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 10980 11354 11008 11630
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10888 11150 10916 11183
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10810 10916 11086
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 10130 10272 10610
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10244 9382 10272 10066
rect 10336 9450 10364 10474
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10336 9194 10364 9386
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10244 9166 10364 9194
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9864 8424 9916 8430
rect 9968 8412 9996 9114
rect 9916 8384 9996 8412
rect 9864 8366 9916 8372
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8772 7342 8800 7958
rect 9692 7342 9720 8366
rect 9876 8022 9904 8366
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 8022 10180 8230
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7546 10180 7958
rect 10244 7886 10272 9166
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8634 10364 8910
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10336 7868 10364 8570
rect 10428 8430 10456 9046
rect 10520 9042 10548 9454
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10612 8022 10640 8774
rect 10704 8634 10732 10406
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 8430 10824 8910
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 8090 10824 8366
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10508 7880 10560 7886
rect 10336 7840 10508 7868
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8772 5234 8800 6054
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8864 5166 8892 6054
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 7484 4758 7512 5102
rect 8864 4826 8892 5102
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 7472 4752 7524 4758
rect 7300 4712 7472 4740
rect 6460 4276 6512 4282
rect 7116 4270 7236 4298
rect 7300 4282 7328 4712
rect 7472 4694 7524 4700
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 6460 4218 6512 4224
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7116 3602 7144 4150
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 5736 3058 5764 3538
rect 6012 3398 6040 3538
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5184 2650 5212 2858
rect 5460 2650 5488 2926
rect 6012 2854 6040 3334
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 7116 2650 7144 3538
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 2410 54 2728 82
rect 4894 60 4950 800
rect 18 0 74 54
rect 2410 0 2466 54
rect 4894 8 4896 60
rect 4948 8 4950 60
rect 7208 82 7236 4270
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7484 4146 7512 4558
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 8128 3126 8156 4694
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 3942 8524 4490
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8588 3398 8616 4626
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3194 8892 3334
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 9232 2990 9260 3946
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3058 9628 3878
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 7576 2650 7604 2926
rect 9784 2922 9812 6190
rect 10152 5914 10180 7278
rect 10244 6934 10272 7822
rect 10336 7342 10364 7840
rect 10508 7822 10560 7828
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10336 6934 10364 7278
rect 10508 6996 10560 7002
rect 10612 6984 10640 7958
rect 10560 6956 10640 6984
rect 10508 6938 10560 6944
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5030 9996 5714
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9876 4282 9904 4626
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10244 3534 10272 6870
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5778 10456 6190
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 11072 5370 11100 9318
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11348 7410 11376 8230
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11716 5778 11744 8230
rect 11900 6934 11928 8842
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11900 6458 11928 6870
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5914 11836 6190
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4282 10916 4966
rect 11152 4684 11204 4690
rect 11256 4672 11284 5578
rect 11716 5370 11744 5714
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 5166 11744 5306
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4690 11376 4966
rect 11204 4644 11284 4672
rect 11152 4626 11204 4632
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3126 10272 3470
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7378 82 7434 800
rect 7208 54 7434 82
rect 4894 0 4950 8
rect 7378 0 7434 54
rect 9862 82 9918 800
rect 10152 82 10180 2790
rect 10244 2650 10272 3062
rect 10612 2650 10640 3606
rect 11256 2990 11284 4644
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11348 3942 11376 4626
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11256 2650 11284 2926
rect 11348 2854 11376 3878
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3194 11560 3606
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11900 2650 11928 3538
rect 12084 3040 12112 11494
rect 12452 11286 12480 11630
rect 12636 11286 12664 12378
rect 12728 12306 12756 13398
rect 12820 13190 12848 13824
rect 12900 13806 12952 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13372 13530 13400 13806
rect 14200 13530 14228 14418
rect 14476 14074 14504 14554
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12820 12170 12848 13126
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 13648 11762 13676 12174
rect 13924 11898 13952 12242
rect 14384 12102 14412 12718
rect 14476 12442 14504 12718
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12636 10810 12664 11222
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9042 12296 9522
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12360 8974 12388 10066
rect 12820 9994 12848 10406
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9586 12940 9862
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8090 12388 8910
rect 12912 8634 12940 9522
rect 13004 9042 13032 9998
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13004 8090 13032 8978
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13096 7993 13124 10542
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13372 9450 13400 9930
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13082 7984 13138 7993
rect 13082 7919 13138 7928
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12360 6390 12388 6870
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6458 12664 6734
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 13004 5778 13032 7142
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13004 5302 13032 5714
rect 13096 5370 13124 5714
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12176 4146 12204 4762
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12084 3012 12204 3040
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11992 2825 12020 2926
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11978 2816 12034 2825
rect 11978 2751 12034 2760
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 9862 54 10180 82
rect 12084 82 12112 2858
rect 12176 1358 12204 3012
rect 12636 2990 12664 4490
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3738 12940 4082
rect 13372 4010 13400 4422
rect 13464 4146 13492 5782
rect 13556 5642 13584 7919
rect 13648 6118 13676 11018
rect 14108 10810 14136 11766
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14108 8974 14136 10746
rect 14752 10266 14780 10746
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14844 9926 14872 15127
rect 15120 14550 15148 16186
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 14936 12714 14964 14486
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 13530 15240 13670
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 11762 14964 12650
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14936 11218 14964 11698
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 15028 9722 15056 9998
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14922 9616 14978 9625
rect 14922 9551 14978 9560
rect 14936 9518 14964 9551
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14660 9042 14688 9386
rect 15028 9178 15056 9658
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14016 6866 14044 8230
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7410 14136 7686
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13556 4758 13584 5578
rect 13648 4826 13676 6054
rect 14108 5778 14136 7346
rect 14844 7342 14872 8230
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14292 6934 14320 7278
rect 14844 7002 14872 7278
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 15028 6322 15056 7142
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5098 14136 5510
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13924 3602 13952 4082
rect 14200 4010 14228 5034
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14292 4078 14320 4490
rect 14568 4146 14596 5102
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14200 3602 14228 3946
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13648 3194 13676 3470
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12636 2650 12664 2926
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12912 2514 12940 3130
rect 13740 2650 13768 3470
rect 14200 2650 14228 3538
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14384 2582 14412 2790
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 12346 82 12402 800
rect 12084 54 12402 82
rect 14568 82 14596 3606
rect 14752 3398 14780 4082
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14936 3738 14964 3946
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14752 2990 14780 3334
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14752 2582 14780 2926
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 15120 1601 15148 11494
rect 15304 10062 15332 19722
rect 15752 19168 15804 19174
rect 15948 19156 15976 19858
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19310 16068 19790
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16132 19174 16160 19722
rect 16776 19514 16804 19858
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16028 19168 16080 19174
rect 15948 19128 16028 19156
rect 15752 19110 15804 19116
rect 16028 19110 16080 19116
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15764 18154 15792 19110
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15948 18290 15976 18770
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15764 17882 15792 18090
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15948 17678 15976 18226
rect 16040 18057 16068 19110
rect 16592 18970 16620 19246
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16026 18048 16082 18057
rect 16026 17983 16082 17992
rect 16408 17678 16436 18702
rect 17328 17746 17356 19178
rect 17788 18970 17816 19858
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17972 18902 18000 19858
rect 18616 19854 18644 20742
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18524 19378 18552 19654
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18248 18630 18276 19246
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 15948 17338 15976 17614
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16408 17066 16436 17614
rect 16500 17338 16528 17682
rect 17328 17338 17356 17682
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17512 17134 17540 17478
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 17512 16726 17540 17070
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15764 16114 15792 16526
rect 16500 16250 16528 16662
rect 17788 16250 17816 17682
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 15162 15884 15438
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15580 13394 15608 13670
rect 15764 13530 15792 14350
rect 15856 14006 15884 15098
rect 15948 14822 15976 15506
rect 17052 14958 17080 15574
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14396 15976 14758
rect 16120 14408 16172 14414
rect 15948 14368 16120 14396
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15856 13394 15884 13942
rect 15948 13938 15976 14368
rect 16120 14350 16172 14356
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16408 13870 16436 14826
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15844 13388 15896 13394
rect 16684 13376 16712 13874
rect 17052 13814 17080 14894
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 16960 13802 17080 13814
rect 16948 13796 17080 13802
rect 17000 13786 17080 13796
rect 16948 13738 17000 13744
rect 16960 13530 16988 13738
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16764 13388 16816 13394
rect 16684 13348 16764 13376
rect 15844 13330 15896 13336
rect 16764 13330 16816 13336
rect 15580 12782 15608 13330
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 12442 15516 12650
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15384 11756 15436 11762
rect 15488 11744 15516 12378
rect 15672 12102 15700 13194
rect 15856 12986 15884 13330
rect 16776 12986 16804 13330
rect 17236 12986 17264 14214
rect 17788 13814 17816 16186
rect 17880 15910 17908 17478
rect 18248 17134 18276 18566
rect 18604 17196 18656 17202
rect 18708 17184 18736 24550
rect 18892 24410 18920 24686
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18892 23730 18920 24346
rect 18984 24274 19012 24686
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 19168 23594 19196 24278
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19168 23322 19196 23530
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 19352 23254 19380 24210
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19996 23322 20024 23666
rect 20364 23662 20392 24142
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 21010 18920 21422
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18892 20602 18920 20946
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19076 18834 19104 19450
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18086 19104 18770
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18656 17156 18736 17184
rect 18604 17138 18656 17144
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18984 17066 19012 17614
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16794 19012 17002
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18248 16046 18276 16730
rect 19076 16658 19104 18022
rect 19168 17882 19196 22442
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19996 22166 20024 23258
rect 20180 23254 20208 23598
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20456 22642 20484 23802
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19260 20942 19288 21422
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19628 20398 19656 20810
rect 20456 20466 20484 20946
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 20364 20330 20392 20402
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 20364 20058 20392 20266
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20456 19990 20484 20402
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19444 19360 19472 19858
rect 19524 19372 19576 19378
rect 19444 19332 19524 19360
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19260 18970 19288 19178
rect 19444 18970 19472 19332
rect 19524 19314 19576 19320
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19444 17882 19472 18294
rect 20456 18222 20484 18702
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18800 15978 18828 16458
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 15162 18460 15506
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18524 14958 18552 15302
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18432 14414 18460 14894
rect 18524 14482 18552 14894
rect 18800 14618 18828 15914
rect 19260 14890 19288 16050
rect 19444 15366 19472 16594
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 20272 15638 20300 17002
rect 20456 16726 20484 18158
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20626 16416 20682 16425
rect 20548 16250 20576 16390
rect 20626 16351 20682 16360
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 20640 15570 20668 16351
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18432 14074 18460 14350
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 17788 13786 17908 13814
rect 18800 13802 18828 14418
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 17880 13394 17908 13786
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17236 12782 17264 12922
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 16316 12442 16344 12718
rect 17236 12442 17264 12718
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15436 11716 15516 11744
rect 15384 11698 15436 11704
rect 15672 11082 15700 12038
rect 15948 11286 15976 12242
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 11626 16068 12038
rect 18248 11762 18276 12718
rect 18432 12306 18460 13330
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16040 11354 16068 11562
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15384 10600 15436 10606
rect 15382 10568 15384 10577
rect 15436 10568 15438 10577
rect 15382 10503 15438 10512
rect 15396 10470 15424 10503
rect 15764 10470 15792 11154
rect 16868 10606 16896 11562
rect 18524 11286 18552 12650
rect 18892 12442 18920 14350
rect 19168 13870 19196 14486
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19168 13530 19196 13806
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19260 13462 19288 13738
rect 19352 13734 19380 14418
rect 19444 14006 19472 15302
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13530 19380 13670
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12714 19012 13126
rect 19260 12850 19288 13398
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11626 19012 12038
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18432 10606 18460 11154
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10606 18552 11018
rect 18616 10742 18644 11562
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15304 9518 15332 9862
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15106 1592 15162 1601
rect 15106 1527 15162 1536
rect 14830 82 14886 800
rect 14568 54 14886 82
rect 15212 66 15240 9318
rect 15304 2854 15332 9454
rect 15580 9382 15608 10066
rect 15764 9926 15792 10406
rect 16868 10130 16896 10542
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17880 10062 17908 10406
rect 18340 10130 18368 10474
rect 18432 10266 18460 10542
rect 18524 10266 18552 10542
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 17420 9722 17448 9998
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15568 9036 15620 9042
rect 15488 8996 15568 9024
rect 15488 8498 15516 8996
rect 15568 8978 15620 8984
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 8401 15516 8434
rect 15474 8392 15530 8401
rect 15474 8327 15530 8336
rect 15764 7954 15792 8774
rect 15856 8430 15884 9386
rect 16684 8974 16712 9454
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8634 16712 8910
rect 16868 8634 16896 9658
rect 17880 9110 17908 9998
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 18156 8498 18184 8978
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 7954 16068 8230
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7410 16988 7890
rect 18156 7750 18184 8434
rect 18248 8430 18276 9386
rect 18340 9178 18368 10066
rect 18432 9722 18460 10202
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18524 9654 18552 10202
rect 19168 10062 19196 10542
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19444 9994 19472 10406
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 19248 8900 19300 8906
rect 19248 8842 19300 8848
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 6798 15976 7142
rect 16316 6798 16344 7346
rect 16960 7002 16988 7346
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15580 6322 15608 6734
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15488 5574 15516 6122
rect 15580 5914 15608 6258
rect 16316 5914 16344 6734
rect 16684 5914 16712 6802
rect 17328 6458 17356 7210
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17788 5914 17816 6870
rect 18156 6798 18184 7686
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 6458 18184 6734
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18248 6322 18276 8366
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18340 6866 18368 7890
rect 18524 7478 18552 8298
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18616 7342 18644 7754
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18616 7002 18644 7278
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18708 6322 18736 7822
rect 18800 7342 18828 8774
rect 19260 8362 19288 8842
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19260 8090 19288 8298
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19444 7954 19472 8774
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7342 19012 7822
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18800 6866 18828 7278
rect 18984 6934 19012 7278
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 18248 5846 18276 6258
rect 18708 5914 18736 6258
rect 19168 6186 19196 6598
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 19168 5914 19196 6122
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5234 15516 5510
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15764 4214 15792 4558
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15856 4078 15884 4966
rect 16132 4078 16160 5034
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4690 16896 4966
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15488 2990 15516 4014
rect 16132 3670 16160 4014
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16316 3602 16344 4558
rect 16868 4282 16896 4626
rect 16960 4486 16988 5782
rect 18248 5166 18276 5782
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 17604 4690 17632 5102
rect 18984 5098 19012 5578
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18984 4826 19012 5034
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19076 4690 19104 5714
rect 19248 5228 19300 5234
rect 19444 5216 19472 7890
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19904 6866 19932 15302
rect 20640 15162 20668 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20272 14482 20300 14826
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19996 13938 20024 14214
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20272 13870 20300 14418
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20088 13734 20116 13806
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20364 10606 20392 11562
rect 20640 11558 20668 12242
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 9722 20576 10542
rect 20640 9722 20668 11494
rect 20732 11257 20760 27254
rect 20810 27171 20866 27254
rect 23124 27254 23350 27282
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22480 24954 22508 25298
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 21192 23866 21220 24210
rect 21468 24070 21496 24686
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 21744 24206 21772 24550
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21192 23254 21220 23530
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22574 21220 22918
rect 21560 22574 21588 22986
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21192 22098 21220 22510
rect 21560 22098 21588 22510
rect 21180 22092 21232 22098
rect 21180 22034 21232 22040
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21100 19922 21128 21286
rect 21192 21146 21220 22034
rect 21560 21554 21588 22034
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21100 19514 21128 19858
rect 21468 19718 21496 20878
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21100 19310 21128 19450
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21376 18426 21404 18702
rect 21468 18630 21496 19654
rect 21744 19174 21772 24142
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 22020 22574 22048 23054
rect 22572 22982 22600 25094
rect 23124 24954 23152 27254
rect 23294 27171 23350 27254
rect 25516 27254 25742 27282
rect 23112 24948 23164 24954
rect 23112 24890 23164 24896
rect 23124 24750 23152 24890
rect 25516 24886 25544 27254
rect 25686 27171 25742 27254
rect 25504 24880 25556 24886
rect 25504 24822 25556 24828
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22664 24313 22692 24346
rect 22650 24304 22706 24313
rect 22650 24239 22706 24248
rect 22664 23866 22692 24239
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22940 23866 22968 24142
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22848 22574 22876 23054
rect 23032 22778 23060 23122
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21836 21078 21864 22374
rect 22020 21146 22048 22510
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21836 20602 21864 21014
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 22112 20262 22140 22102
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 21486 22232 21830
rect 22848 21690 22876 22510
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22848 21486 22876 21626
rect 23032 21554 23060 22714
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21914 20088 21970 20097
rect 21914 20023 21970 20032
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20916 17202 20944 17818
rect 21468 17678 21496 18566
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 14958 20944 15914
rect 21008 15706 21036 17478
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21100 16726 21128 17070
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21192 16454 21220 17070
rect 21468 16998 21496 17614
rect 21744 17270 21772 17614
rect 21836 17542 21864 18838
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16182 21220 16390
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21928 15570 21956 20023
rect 22204 19922 22232 21422
rect 22572 21146 22600 21422
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22388 20602 22416 21014
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22388 19514 22416 20538
rect 22572 19990 22600 21082
rect 23032 20942 23060 21490
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22756 19514 22784 19858
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 18222 22324 19246
rect 22756 18902 22784 19450
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22480 17814 22508 18022
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22296 16046 22324 16594
rect 22388 16590 22416 17614
rect 22480 17338 22508 17750
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22664 16658 22692 17070
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22388 16114 22416 16526
rect 22572 16182 22600 16526
rect 22664 16250 22692 16594
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22388 15570 22416 16050
rect 22572 15638 22600 16118
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20916 14278 20944 14894
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 21376 14006 21404 14350
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 20916 11354 20944 13942
rect 21376 13814 21404 13942
rect 21100 13786 21404 13814
rect 21100 12306 21128 13786
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20718 11248 20774 11257
rect 20718 11183 20774 11192
rect 21100 11082 21128 12242
rect 21376 11694 21404 13398
rect 21468 12782 21496 15302
rect 21928 15162 21956 15506
rect 22388 15162 22416 15506
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22204 14550 22232 14758
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 13734 22140 14350
rect 22204 14074 22232 14486
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13462 22140 13670
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21560 12646 21588 13330
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21744 12374 21772 12582
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 11830 21680 12174
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21744 11694 21772 12310
rect 22020 11694 22048 12650
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 21376 11218 21404 11630
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21088 11076 21140 11082
rect 21140 11036 21220 11064
rect 21088 11018 21140 11024
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20180 7993 20208 9454
rect 21100 9382 21128 10066
rect 21192 9450 21220 11036
rect 21284 10470 21312 11154
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 9518 21312 10406
rect 21376 10266 21404 11154
rect 22020 11082 22048 11630
rect 22112 11354 22140 12310
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 22020 10266 22048 11018
rect 22112 10810 22140 11290
rect 22204 11286 22232 11630
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22388 10674 22416 14894
rect 22940 14006 22968 16934
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23400 14550 23428 15846
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 25042 13288 25098 13297
rect 25042 13223 25098 13232
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 22480 11218 22508 12718
rect 23400 12374 23428 12718
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 22480 10810 22508 11154
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8634 21128 9318
rect 21192 8974 21220 9386
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21744 8294 21772 8910
rect 21836 8498 21864 9318
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 20166 7984 20222 7993
rect 20166 7919 20222 7928
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20456 7546 20484 7890
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5846 19932 6802
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19524 5228 19576 5234
rect 19444 5188 19524 5216
rect 19248 5170 19300 5176
rect 19524 5170 19576 5176
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16960 3602 16988 4422
rect 17604 4282 17632 4626
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17972 4078 18000 4422
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16316 3194 16344 3538
rect 16960 3194 16988 3538
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17236 3058 17264 3470
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15488 2650 15516 2926
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 17314 82 17370 800
rect 17420 82 17448 3878
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17696 3194 17724 3606
rect 19076 3602 19104 4626
rect 19260 4010 19288 5170
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19996 4758 20024 6598
rect 20824 6322 20852 7278
rect 21560 6934 21588 7278
rect 21744 7274 21772 8230
rect 22296 8090 22324 9046
rect 22388 8090 22416 10610
rect 22664 10520 22692 11154
rect 23032 10810 23060 11154
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22744 10532 22796 10538
rect 22664 10492 22744 10520
rect 22664 10130 22692 10492
rect 22744 10474 22796 10480
rect 23032 10266 23060 10746
rect 25056 10577 25084 13223
rect 25042 10568 25098 10577
rect 25042 10503 25098 10512
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22664 9722 22692 10066
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22756 8294 22784 8774
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20456 5778 20484 6122
rect 20824 5914 20852 6258
rect 21100 6186 21128 6734
rect 21560 6254 21588 6870
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6458 21864 6734
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 22020 6236 22048 6598
rect 22100 6248 22152 6254
rect 22020 6208 22100 6236
rect 21088 6180 21140 6186
rect 21088 6122 21140 6128
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20824 4826 20852 5850
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17696 2650 17724 3130
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 18984 2446 19012 3470
rect 19076 2650 19104 3538
rect 19444 3058 19472 4626
rect 19628 4078 19656 4694
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 19996 4146 20024 4422
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19996 3398 20024 4082
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 9862 0 9918 54
rect 12346 0 12402 54
rect 14830 0 14886 54
rect 15200 60 15252 66
rect 15200 2 15252 8
rect 17314 54 17448 82
rect 19798 82 19854 800
rect 19904 82 19932 2858
rect 19996 2650 20024 3334
rect 20364 3194 20392 4014
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20456 2990 20484 3878
rect 20640 2990 20668 4422
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20916 3534 20944 3946
rect 21100 3534 21128 6122
rect 21560 5914 21588 6190
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 22020 5846 22048 6208
rect 22100 6190 22152 6196
rect 22756 6186 22784 8230
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22940 6458 22968 6802
rect 23124 6497 23152 9318
rect 23400 9110 23428 9658
rect 25042 9616 25098 9625
rect 25042 9551 25098 9560
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 25056 8401 25084 9551
rect 25042 8392 25098 8401
rect 24492 8356 24544 8362
rect 25042 8327 25098 8336
rect 24492 8298 24544 8304
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 7546 23244 7890
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23110 6488 23166 6497
rect 22928 6452 22980 6458
rect 23308 6458 23336 7686
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23110 6423 23166 6432
rect 23296 6452 23348 6458
rect 22928 6394 22980 6400
rect 23296 6394 23348 6400
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21468 5370 21496 5578
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21836 5166 21864 5714
rect 22020 5370 22048 5782
rect 22848 5778 22876 6190
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22848 5574 22876 5714
rect 23584 5642 23612 6734
rect 23572 5636 23624 5642
rect 23572 5578 23624 5584
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21836 4826 21864 5102
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 22848 4758 22876 5510
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 23584 4690 23612 5578
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4078 21680 4558
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21928 4146 21956 4422
rect 22480 4282 22508 4626
rect 23584 4282 23612 4626
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21468 3534 21496 4014
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20640 2650 20668 2926
rect 21100 2922 21128 3470
rect 21376 3126 21404 3470
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 21376 2650 21404 3062
rect 21468 2650 21496 3470
rect 21836 3194 21864 3606
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22020 2990 22048 4014
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3194 22692 3878
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 22376 1352 22428 1358
rect 22376 1294 22428 1300
rect 19798 54 19932 82
rect 22282 82 22338 800
rect 22388 82 22416 1294
rect 22282 54 22416 82
rect 24504 82 24532 8298
rect 24766 82 24822 800
rect 24504 54 24822 82
rect 17314 0 17370 54
rect 19798 0 19854 54
rect 22282 0 22338 54
rect 24766 0 24822 54
<< via2 >>
rect 1674 25064 1730 25120
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 1214 21392 1270 21448
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 1214 9560 1270 9616
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 1674 10376 1730 10432
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 1582 7792 1638 7848
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 10414 15000 10470 15056
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 12070 15136 12126 15192
rect 14830 15136 14886 15192
rect 10874 11192 10930 11248
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 13082 7928 13138 7984
rect 13542 7928 13598 7984
rect 11978 2760 12034 2816
rect 14922 9560 14978 9616
rect 16026 17992 16082 18048
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 20626 16360 20682 16416
rect 15382 10548 15384 10568
rect 15384 10548 15436 10568
rect 15436 10548 15438 10568
rect 15382 10512 15438 10548
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 15106 1536 15162 1592
rect 15474 8336 15530 8392
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 22650 24248 22706 24304
rect 21914 20032 21970 20088
rect 20718 11192 20774 11248
rect 25042 13232 25098 13288
rect 20166 7928 20222 7984
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 25042 10512 25098 10568
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 25042 9560 25098 9616
rect 25042 8336 25098 8392
rect 23110 6432 23166 6488
<< metal3 >>
rect 0 25576 800 25696
rect 19568 25600 19888 25601
rect 62 25122 122 25576
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 1669 25122 1735 25125
rect 62 25120 1735 25122
rect 62 25064 1674 25120
rect 1730 25064 1735 25120
rect 62 25062 1735 25064
rect 1669 25059 1735 25062
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 22645 24306 22711 24309
rect 25027 24306 25827 24336
rect 22645 24304 25827 24306
rect 22645 24248 22650 24304
rect 22706 24248 25827 24304
rect 22645 24246 25827 24248
rect 22645 24243 22711 24246
rect 25027 24216 25827 24246
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 0 21904 800 22024
rect 62 21450 122 21904
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 1209 21450 1275 21453
rect 62 21448 1275 21450
rect 62 21392 1214 21448
rect 1270 21392 1275 21448
rect 62 21390 1275 21392
rect 1209 21387 1275 21390
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 25027 20544 25827 20664
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 21909 20090 21975 20093
rect 25086 20090 25146 20544
rect 21909 20088 25146 20090
rect 21909 20032 21914 20088
rect 21970 20032 25146 20088
rect 21909 20030 25146 20032
rect 21909 20027 21975 20030
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 0 18232 800 18352
rect 62 18050 122 18232
rect 16021 18050 16087 18053
rect 62 18048 16087 18050
rect 62 17992 16026 18048
rect 16082 17992 16087 18048
rect 62 17990 16087 17992
rect 16021 17987 16087 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 25027 16872 25827 16992
rect 19568 16831 19888 16832
rect 20621 16418 20687 16421
rect 25086 16418 25146 16872
rect 20621 16416 25146 16418
rect 20621 16360 20626 16416
rect 20682 16360 25146 16416
rect 20621 16358 25146 16360
rect 20621 16355 20687 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 12065 15194 12131 15197
rect 14825 15194 14891 15197
rect 12065 15192 14891 15194
rect 12065 15136 12070 15192
rect 12126 15136 14830 15192
rect 14886 15136 14891 15192
rect 12065 15134 14891 15136
rect 12065 15131 12131 15134
rect 14825 15131 14891 15134
rect 10409 15058 10475 15061
rect 62 15056 10475 15058
rect 62 15000 10414 15056
rect 10470 15000 10475 15056
rect 62 14998 10475 15000
rect 62 14680 122 14998
rect 10409 14995 10475 14998
rect 19568 14720 19888 14721
rect 0 14560 800 14680
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 25027 13290 25827 13320
rect 24956 13288 25827 13290
rect 24956 13232 25042 13288
rect 25098 13232 25827 13288
rect 24956 13230 25827 13232
rect 25027 13200 25827 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 10869 11250 10935 11253
rect 20713 11250 20779 11253
rect 10869 11248 20779 11250
rect 10869 11192 10874 11248
rect 10930 11192 20718 11248
rect 20774 11192 20779 11248
rect 10869 11190 20779 11192
rect 10869 11187 10935 11190
rect 20713 11187 20779 11190
rect 0 10888 800 11008
rect 4208 10912 4528 10913
rect 62 10434 122 10888
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 15377 10570 15443 10573
rect 25037 10570 25103 10573
rect 15377 10568 25103 10570
rect 15377 10512 15382 10568
rect 15438 10512 25042 10568
rect 25098 10512 25103 10568
rect 15377 10510 25103 10512
rect 15377 10507 15443 10510
rect 25037 10507 25103 10510
rect 1669 10434 1735 10437
rect 62 10432 1735 10434
rect 62 10376 1674 10432
rect 1730 10376 1735 10432
rect 62 10374 1735 10376
rect 1669 10371 1735 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 1209 9618 1275 9621
rect 14917 9618 14983 9621
rect 25027 9618 25827 9648
rect 1209 9616 14983 9618
rect 1209 9560 1214 9616
rect 1270 9560 14922 9616
rect 14978 9560 14983 9616
rect 1209 9558 14983 9560
rect 24956 9616 25827 9618
rect 24956 9560 25042 9616
rect 25098 9560 25827 9616
rect 24956 9558 25827 9560
rect 1209 9555 1275 9558
rect 14917 9555 14983 9558
rect 25027 9528 25827 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 15469 8394 15535 8397
rect 25037 8394 25103 8397
rect 15469 8392 25103 8394
rect 15469 8336 15474 8392
rect 15530 8336 25042 8392
rect 25098 8336 25103 8392
rect 15469 8334 25103 8336
rect 15469 8331 15535 8334
rect 25037 8331 25103 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 13077 7986 13143 7989
rect 13537 7986 13603 7989
rect 20161 7986 20227 7989
rect 13077 7984 20227 7986
rect 13077 7928 13082 7984
rect 13138 7928 13542 7984
rect 13598 7928 20166 7984
rect 20222 7928 20227 7984
rect 13077 7926 20227 7928
rect 13077 7923 13143 7926
rect 13537 7923 13603 7926
rect 20161 7923 20227 7926
rect 1577 7850 1643 7853
rect 62 7848 1643 7850
rect 62 7792 1582 7848
rect 1638 7792 1643 7848
rect 62 7790 1643 7792
rect 62 7336 122 7790
rect 1577 7787 1643 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 0 7216 800 7336
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 23105 6490 23171 6493
rect 23105 6488 25146 6490
rect 23105 6432 23110 6488
rect 23166 6432 25146 6488
rect 23105 6430 25146 6432
rect 23105 6427 23171 6430
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 25086 5976 25146 6430
rect 19568 5951 19888 5952
rect 25027 5856 25827 5976
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3544 800 3664
rect 62 2818 122 3544
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 11973 2818 12039 2821
rect 62 2816 12039 2818
rect 62 2760 11978 2816
rect 12034 2760 12039 2816
rect 62 2758 12039 2760
rect 11973 2755 12039 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 25027 2184 25827 2304
rect 4208 2143 4528 2144
rect 15101 1594 15167 1597
rect 25086 1594 25146 2184
rect 15101 1592 25146 1594
rect 15101 1536 15106 1592
rect 15162 1536 25146 1592
rect 15101 1534 25146 1536
rect 15101 1531 15167 1534
<< via3 >>
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
<< metal4 >>
rect 4208 25056 4528 25616
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5576 4528 6496
rect 4208 5472 4250 5576
rect 4486 5472 4528 5576
rect 4208 5408 4216 5472
rect 4520 5408 4528 5472
rect 4208 5340 4250 5408
rect 4486 5340 4528 5408
rect 4208 4384 4528 5340
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 25600 19888 25616
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20894 19888 21184
rect 19568 20658 19610 20894
rect 19846 20658 19888 20894
rect 19568 20160 19888 20658
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
<< via4 >>
rect 4250 5472 4486 5576
rect 4250 5408 4280 5472
rect 4280 5408 4296 5472
rect 4296 5408 4360 5472
rect 4360 5408 4376 5472
rect 4376 5408 4440 5472
rect 4440 5408 4456 5472
rect 4456 5408 4486 5472
rect 4250 5340 4486 5408
rect 19610 20658 19846 20894
<< metal5 >>
rect 1104 20894 24656 20936
rect 1104 20658 19610 20894
rect 19846 20658 24656 20894
rect 1104 20616 24656 20658
rect 1104 5576 24656 5618
rect 1104 5340 4250 5576
rect 4486 5340 24656 5576
rect 1104 5298 24656 5340
use scs8hd_fill_2  FILLER_1_8 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_3 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_9 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__430__A /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__430__B
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_and2_4  _430_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 682 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_17 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__351__A
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_12 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_29
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_24
timestamp 1586364061
transform 1 0 3312 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__431__A
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _351_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__B1
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__A2
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__432__A1
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _431_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_45
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__A
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _427_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__434__A
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_61
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__426__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__434__B
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _426_
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use scs8hd_decap_12  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_77 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__633__CLK
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__447__A
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_and2_4  _447_
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 682 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__634__CLK
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_103
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_105
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__634__D
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__634__RESETB
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__447__B
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_112
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__424__A
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _424_
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__B2
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__338__B
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_120
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__339__A
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _339_
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 314 592
use scs8hd_and2_4  _338_
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 682 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__A2
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__A1
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__338__A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__B1
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_xor2_4  _342_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 2062 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__342__B
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__342__A
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__336__A
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__694__CLK
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__694__RESETB
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__694__D
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__632__A
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_184
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__619__A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _353_
timestamp 1586364061
transform 1 0 18492 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_200
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__353__A
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__619__B
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _632_
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_and2_4  _619_
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 682 592
use scs8hd_decap_4  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__A1N
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_a2bb2o_4  _334_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_1_224
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__631__A
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__691__D
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_228
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__B2
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__B1
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__691__RESETB
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _631_
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__691__CLK
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_245
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 24656 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 24656 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__638__RESETB
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__432__B2
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_o22a_4  _432_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__433__B1
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_xor2_4  _434_
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 2062 592
use scs8hd_decap_6  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_85
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__448__A
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_dfrtp_4  _634_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__696__D
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_o22a_4  _340_
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 1326 592
use scs8hd_decap_6  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__341__A2N
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _336_
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_1  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use scs8hd_dfrtp_4  _694_
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__334__A2N
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__356__A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_1  _356_
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_dfrtp_4  _691_
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_2_252
timestamp 1586364061
transform 1 0 24288 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 24656 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__638__D
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_dfrtp_4  _638_
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__433__A2N
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__433__A1N
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__633__RESETB
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_dfrtp_4  _633_
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__425__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__468__A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__604__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__468__B
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_and2_4  _468_
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 682 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_dfrtp_4  _696_
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__693__D
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_a2bb2o_4  _341_
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__355__A
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__693__RESETB
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_xor2_4  _335_
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__333__B1
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__620__A
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__617__A
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_o22a_4  _333_
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 1326 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 24656 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__444__B
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__444__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__443__B2
timestamp 1586364061
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__638__CLK
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__439__A
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_37
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _420_
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__420__A
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__433__B2
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_70
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__633__D
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_a2bb2o_4  _433_
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__639__CLK
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__639__RESETB
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_1  _448_
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_1  _425_
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_98
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_1  _604_
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_120
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__696__CLK
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__A
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__696__RESETB
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _350_
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_151
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__693__CLK
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__341__B1
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_dfrtp_4  _693_
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__335__B
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _355_
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__A
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__357__A
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__333__A2
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__A1
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_221
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__621__A1
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _620_
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_233
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_225
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__B2
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__621__B2
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _617_
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 24656 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_xor2_4  _444_
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__640__D
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__640__RESETB
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__640__CLK
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__450__B2
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__450__B1
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__450__A2N
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__450__A1N
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__639__D
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_dfrtp_4  _639_
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__469__A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__A
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__428__A
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _428_
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__349__A
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _352_
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__A
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__349__B
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__337__A
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__341__B2
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__341__A1N
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _337_
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 866 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_181
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_172
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__354__A
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__692__D
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_dfrtp_4  _692_
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 2154 592
use scs8hd_buf_1  _354_
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_209
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 590 592
use scs8hd_decap_6  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_222
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__618__A
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__621__A2
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__621__B1
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _618_
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 24656 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__443__A1N
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__637__RESETB
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_8
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__443__A2N
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__637__D
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_8  _439_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_dfrtp_4  _637_
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_37
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__637__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__451__A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_dfrtp_4  _640_
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 2154 592
use scs8hd_buf_1  _418_
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_57
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__A2
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__418__A
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__B1
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_a2bb2o_4  _450_
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 1510 592
use scs8hd_o22a_4  _449_
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__445__A
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__449__B2
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__419__A
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _419_
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__A
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__636__RESETB
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _469_
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _416_
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__A
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__636__D
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _422_
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_buf_1  _358_
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_99
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__695__CLK
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__636__CLK
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_xor2_4  _349_
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__695__RESETB
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__695__D
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__A1
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__B1
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_dfrtp_4  _695_
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_170
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__628__B2
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__690__CLK
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__692__CLK
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__628__A1
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__628__A2
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__628__B1
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__692__RESETB
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__690__D
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 406 592
use scs8hd_dfrtp_4  _690_
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_6_194
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _357_
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_198
timestamp 1586364061
transform 1 0 19320 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__332__A
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__622__B1
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_212
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_221
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__622__A1N
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__687__D
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_237
timestamp 1586364061
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__687__RESETB
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_a2bb2o_4  _622_
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1510 592
use scs8hd_o22a_4  _621_
timestamp 1586364061
transform 1 0 21620 0 -1 5984
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__687__CLK
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__622__B2
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 24656 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 24656 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_21
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__443__B1
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_a2bb2o_4  _443_
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_8_38
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_25
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__B2
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__451__B
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_xor2_4  _451_
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__449__A1
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _445_
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__645__RESETB
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__645__CLK
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__466__A
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_dfrtp_4  _636_
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__348__A2N
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__B2
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__A2
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_o22a_4  _347_
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__630__A
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__629__A2N
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_o22a_4  _628_
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__623__B
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__690__RESETB
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _332_
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_220
timestamp 1586364061
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__622__A2N
timestamp 1586364061
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use scs8hd_dfrtp_4  _687_
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 2154 592
use scs8hd_decap_8  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 24656 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__B1
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_o22a_4  _442_
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 1326 592
use scs8hd_decap_12  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__417__A
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__421__A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__438__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _421_
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_67
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__446__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__472__A
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__411__A
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_xor2_4  _472_
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 2062 592
use scs8hd_decap_8  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use scs8hd_decap_4  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__645__D
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _466_
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_9_139
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__348__B2
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__348__A1N
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_a2bb2o_4  _348_
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__343__A
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _343_
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__629__A1N
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_a2bb2o_4  _629_
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_202
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__623__A
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__360__A
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_xor2_4  _623_
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__362__A
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 24656 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_11
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__A1
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__440__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_8  _438_
timestamp 1586364061
transform 1 0 2300 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_6  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_6  FILLER_10_37
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__641__CLK
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__415__A
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_1  _417_
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__460__A
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__646__RESETB
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _446_
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__472__B
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__A
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _411_
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__470__A1
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_dfrtp_4  _645_
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_10_118
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__437__A1
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__348__B1
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__437__A2
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_159
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__A
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__630__B
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_1  _346_
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_xor2_4  _630_
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__629__B2
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__624__A
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _625_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_231
timestamp 1586364061
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__A
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__688__RESETB
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _361_
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _360_
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 24656 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _362_
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_8
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _441_
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__442__A2
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__440__B
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__642__RESETB
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__642__D
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_dfrtp_4  _642_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__646__D
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_dfrtp_4  _646_
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__B1
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_a2bb2o_4  _471_
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 1510 592
use scs8hd_fill_1  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__A1N
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__373__A
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_128
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_buf_1  _373_
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__437__B1N
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__344__A
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _344_
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__345__A
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__345__B
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _627_
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__629__B1
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__627__A
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__689__D
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_dfrtp_4  _689_
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__569__A
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__688__CLK
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__688__D
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__569__B
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_and2_4  _569_
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 682 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 24656 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__457__A2N
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__641__RESETB
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_and2_4  _440_
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 682 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__457__B1
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__642__CLK
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__452__A
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  _415_
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__464__B2
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__463__A2
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__463__A1
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _460_
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__646__CLK
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _412_
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__471__A2N
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_o22a_4  _470_
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 1326 592
use scs8hd_decap_8  FILLER_12_113
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_109
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__A2
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 1142 592
use scs8hd_a21boi_4  _437_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 1418 592
use scs8hd_decap_6  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__576__A
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_and2_4  _345_
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 682 592
use scs8hd_fill_1  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__571__A1
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__561__A
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__571__A2
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__689__RESETB
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _624_
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__625__A
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use scs8hd_dfrtp_4  _688_
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 24656 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__457__A1N
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__441__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__641__D
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_dfrtp_4  _641_
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 2154 592
use scs8hd_a2bb2o_4  _457_
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__457__B2
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 406 592
use scs8hd_inv_8  _452_
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__464__B1
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__465__A
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__456__B2
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__464__A2N
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__464__A1N
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__463__B1
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_a2bb2o_4  _464_
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 1510 592
use scs8hd_o22a_4  _463_
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_78
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__414__A
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__459__A
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _414_
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__463__B2
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__B1
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _467_
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__471__B2
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__470__B2
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__429__A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _429_
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__436__A
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__467__A
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__635__CLK
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__635__D
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__635__RESETB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_or2_4  _436_ /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 682 592
use scs8hd_decap_8  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__436__B
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_dfrtp_4  _635_
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__626__A
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__626__B
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_151
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_and2_4  _626_
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 682 592
use scs8hd_and2_4  _576_
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 682 592
use scs8hd_decap_4  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__576__B
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_174
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_170
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__571__B2
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__573__A
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__571__B1
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _561_
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__572__B2
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__572__B1
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_o22a_4  _571_
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 1326 592
use scs8hd_decap_8  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_192
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__689__CLK
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__572__A2N
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__359__A
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _359_
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_220
timestamp 1586364061
transform 1 0 21344 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__615__B2
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__570__A
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _570_
timestamp 1586364061
transform 1 0 21068 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_229
timestamp 1586364061
transform 1 0 22172 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__614__A1
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__562__A
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _611_
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 866 592
use scs8hd_and2_4  _562_
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 682 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__562__B
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_250
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_242
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__611__A
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 24656 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 24656 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_xor2_4  _458_
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__456__B1
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_o22a_4  _456_
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__465__B
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__456__A2
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__643__D
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_dfrtp_4  _643_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__475__A
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _409_
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__CTS_buf_1_0_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__A
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__CTS_root_A
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_clkbuf_4  _CTS_buf_1_0 /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_128
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _423_
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__423__A
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__CTS_buf_1_48_A
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__435__A
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__568__A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__577__A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__435__B
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _568_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_and2_4  _435_
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__572__A1N
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_a2bb2o_4  _572_
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__567__A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _567_
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__366__A
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _364_
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__614__B1
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__614__A2
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__364__A
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_249
timestamp 1586364061
transform 1 0 24012 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__614__B2
timestamp 1586364061
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 24656 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _455_
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_8
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__A
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__455__A
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__458__A
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_20
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__458__B
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_24
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__456__A1
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__644__RESETB
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_xor2_4  _465_
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__643__RESETB
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _459_
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  _475_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_98
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__511__A
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_clkbuf_16  _CTS_root /openLANE_flow/pdks//EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1878 592
use scs8hd_decap_6  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_8  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 774 592
use scs8hd_clkbuf_4  _CTS_buf_1_48
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__676__CLK
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__676__RESETB
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  _577_
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__376__A
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__573__B
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use scs8hd_xor2_4  _573_
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__685__CLK
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__615__A2N
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__685__RESETB
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use scs8hd_o22a_4  _614_
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1326 592
use scs8hd_buf_1  _366_
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 24656 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__644__D
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__454__B
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_inv_8  _453_
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 866 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_dfrtp_4  _644_
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 2154 592
use scs8hd_decap_6  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__643__CLK
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__512__A
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__462__A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _462_
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__461__A
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_and2_4  _461_
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 682 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__461__B
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__511__B
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_and2_4  _511_
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 682 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_128
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__518__A
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_and2_4  _519_
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 682 592
use scs8hd_buf_1  _518_
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__519__B
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_dfrtp_4  _676_
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__673__D
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_dfrtp_4  _673_
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__563__A
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__615__A1N
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__685__D
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_a2bb2o_4  _615_
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1510 592
use scs8hd_decap_4  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__615__B1
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 24656 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_16
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__453__A
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__506__B2
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__506__A2
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_and2_4  _454_
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 682 592
use scs8hd_fill_2  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_24
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__644__CLK
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__413__A
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_1  _413_
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__514__A2N
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__509__A
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_90
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_1  _512_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_99
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__523__A
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_xor2_4  _523_
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__CTS_buf_1_16_A
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__520__A
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__519__A
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _520_
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__580__B
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__B1
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__676__D
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _376_
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__B2
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_179
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__673__CLK
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__A
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__673__RESETB
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__616__A
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__A
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_1  _563_
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_1  _379_
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use scs8hd_dfrtp_4  _685_
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_243
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 24656 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__B
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_and2_4  _504_
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 682 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__504__A
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__506__B1
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _503_
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_20
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_20
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__658__CLK
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__658__RESETB
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_28
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_24
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__503__A
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__505__A
timestamp 1586364061
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__515__A
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__515__B
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _410_
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 314 592
use scs8hd_xor2_4  _515_
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__A1N
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__410__A
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__657__RESETB
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_inv_8  _509_
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use scs8hd_a2bb2o_4  _514_
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 1510 592
use scs8hd_decap_6  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_76
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__B2
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__514__B1
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__510__A
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_90
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__660__CLK
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__660__D
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_dfrtp_4  _660_
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__CTS_buf_1_32_A
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__523__B
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__660__RESETB
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_clkbuf_4  _CTS_buf_1_16
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__A2N
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__B2
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__B1
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 590 592
use scs8hd_clkbuf_4  _CTS_buf_1_32
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__580__A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__377__A
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_xor2_4  _580_
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_151
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__A2
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__A1N
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_a2bb2o_4  _579_
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1510 592
use scs8hd_decap_4  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_172
timestamp 1586364061
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__B2
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__674__CLK
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__579__A2N
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_181
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__564__B2
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__674__RESETB
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__674__D
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  _378_
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 314 592
use scs8hd_dfrtp_4  _674_
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__564__A1
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__565__A2N
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__564__A2
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_209
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__616__B
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__613__A
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__610__A
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_xor2_4  _616_
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 2062 592
use scs8hd_buf_1  _613_
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 314 592
use scs8hd_inv_8  _610_
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 24656 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 24656 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_8
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__658__D
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_dfrtp_4  _658_
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 2154 592
use scs8hd_buf_1  _505_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__502__A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__513__B1
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__657__D
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_dfrtp_4  _657_
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 2154 592
use scs8hd_buf_1  _397_
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__513__B2
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _510_
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__522__A1N
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__A
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__659__RESETB
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__659__D
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_a2bb2o_4  _522_
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_146
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__675__RESETB
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__B1
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__675__D
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_o22a_4  _578_
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__565__B2
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_181
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__565__B1
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_189
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__565__A1N
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__686__RESETB
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__564__B1
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_o22a_4  _564_
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 1326 592
use scs8hd_decap_6  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_234
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__560__A
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__686__CLK
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__686__D
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _560_
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 24656 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__655__RESETB
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_o22a_4  _506_
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 1326 592
use scs8hd_fill_1  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__506__A1
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _502_
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__657__CLK
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__513__A1
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__397__A
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_o22a_4  _513_
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_77
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__526__A
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__659__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_dfrtp_4  _659_
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 2154 592
use scs8hd_buf_1  _396_
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_22_131
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__516__A
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _377_
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_151
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__675__CLK
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_dfrtp_4  _675_
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__566__A
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_a2bb2o_4  _565_
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__559__A
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use scs8hd_dfrtp_4  _686_
timestamp 1586364061
transform 1 0 21344 0 -1 14688
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_243
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 24656 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__655__D
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_dfrtp_4  _655_
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_23_46
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__647__D
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _400_
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__647__RESETB
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__A
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__647__CLK
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__513__A2
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _398_
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_72
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__398__A
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__526__B
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_and2_4  _526_
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 682 592
use scs8hd_fill_2  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__521__A2
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__A
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__B1
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__521__B2
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_o22a_4  _521_
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__578__A1
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__574__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _575_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_inv_8  _517_
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__365__A
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_xor2_4  _566_
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_23_212
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__331__B
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _559_
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__602__A
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__612__B
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _363_
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__363__A
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 24656 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__A2N
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_a2bb2o_4  _507_
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_25
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__B1
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__479__B1
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_dfrtp_4  _647_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__648__CLK
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__648__D
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_72
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__395__A
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__554__A
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__662__D
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _394_
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_137
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__521__A1
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _516_
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_6  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__517__A
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _574_
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_181
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_173
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__575__A
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__566__B
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _365_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__331__A
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__A
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_and2_4  _331_
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 682 592
use scs8hd_decap_4  FILLER_24_229
timestamp 1586364061
transform 1 0 22172 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_225
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__612__A
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use scs8hd_and2_4  _612_
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 682 592
use scs8hd_inv_8  _602_
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  FILLER_24_250
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 24656 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_xor2_4  _508_
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_25_37
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__479__A2N
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__B1
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_o22a_4  _478_
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__479__A1N
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_dfrtp_4  _648_
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_89
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__388__A
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__662__CLK
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__662__RESETB
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__554__B
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_and2_4  _554_
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 682 592
use scs8hd_fill_1  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_128
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__555__A
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_buf_1  _555_
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 314 592
use scs8hd_buf_1  _374_
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__A
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__672__CLK
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_157
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__672__D
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__672__RESETB
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _380_
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_181
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__380__A
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__671__RESETB
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_dfrtp_4  _671_
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_209
timestamp 1586364061
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__603__A
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__B2
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__A2
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__A1
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__607__B1
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _603_
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 24656 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_9
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__507__A1N
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__650__RESETB
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__650__D
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_21
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_17
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_13
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__655__CLK
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__508__B
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__508__A
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_dfrtp_4  _650_
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_25
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__474__A
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__A2
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_38
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_37
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__478__A1
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__399__A
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _474_
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 866 592
use scs8hd_a2bb2o_4  _479_
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__480__A
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__473__A
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__479__B2
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__648__RESETB
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_8  _473_
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_82
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__402__A
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _395_
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_87
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__530__A
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__527__A
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _388_
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 314 592
use scs8hd_xor2_4  _530_
timestamp 1586364061
transform 1 0 9292 0 1 16864
box -38 -48 2062 592
use scs8hd_decap_3  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_98
timestamp 1586364061
transform 1 0 10120 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__605__A
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__A
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_dfrtp_4  _662_
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__381__A
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _381_
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_134
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__557__B2
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__557__B1
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__557__A1N
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__605__B
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_a2bb2o_4  _557_
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_151
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_148
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__556__A1
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__556__B1
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _553_
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 866 592
use scs8hd_dfrtp_4  _672_
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__382__A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_181
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__671__CLK
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__678__D
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__671__D
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__678__CLK
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_dfrtp_4  _678_
timestamp 1586364061
transform 1 0 18216 0 1 16864
box -38 -48 2154 592
use scs8hd_decap_8  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_192
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _372_
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_208
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__608__B2
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_213
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_209
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__608__A2N
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__683__D
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__608__A1N
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__683__CLK
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__683__RESETB
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_237
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use scs8hd_a2bb2o_4  _608_
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 1510 592
use scs8hd_o22a_4  _607_
timestamp 1586364061
transform 1 0 21620 0 -1 16864
box -38 -48 1326 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_249
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 24656 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 24656 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__507__B2
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_14
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__656__RESETB
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__656__CLK
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__406__A
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__650__CLK
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_37
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _399_
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__478__B2
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__480__B
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_48
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use scs8hd_xor2_4  _480_
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__403__A
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _402_
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__530__B
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_1  _527_
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_116
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_98
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__661__CLK
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__529__B1
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__661__RESETB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _392_
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_140
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__557__A2N
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use scs8hd_and2_4  _605_
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 682 592
use scs8hd_fill_2  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__556__A2
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__669__RESETB
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_o22a_4  _556_
timestamp 1586364061
transform 1 0 15456 0 -1 17952
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_174
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_170
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__553__A
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__556__B2
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__678__RESETB
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _382_
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_195
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_191
timestamp 1586364061
transform 1 0 18676 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__375__A
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_1  _375_
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_203
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_28_199
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__609__A
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_209
timestamp 1586364061
transform 1 0 20332 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__608__B1
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__684__RESETB
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use scs8hd_dfrtp_4  _683_
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_244
timestamp 1586364061
transform 1 0 23552 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 24656 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__656__D
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_dfrtp_4  _656_
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__496__A
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__B2
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__A1N
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_52
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_48
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__500__A2N
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__500__B1
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_67
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _401_
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__A
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__529__B2
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__408__A
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _408_
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_89
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__529__A2N
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__529__A1N
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_a2bb2o_4  _529_
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 1510 592
use scs8hd_decap_6  FILLER_29_115
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__661__D
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__669__D
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_dfrtp_4  _669_
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_29_189
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__552__A
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _606_
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__606__A
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__371__A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_xor2_4  _609_
timestamp 1586364061
transform 1 0 19504 0 1 17952
box -38 -48 2062 592
use scs8hd_decap_6  FILLER_29_237
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_233
timestamp 1586364061
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_222
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__A
timestamp 1586364061
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__684__D
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _367_
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_243
timestamp 1586364061
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 24656 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__A2N
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_16
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__487__A
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__481__A
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_buf_1  _406_
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_37
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__499__A2
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__A1
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_a2bb2o_4  _500_
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 1510 592
use scs8hd_decap_4  FILLER_30_66
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__495__A
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_1  _403_
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_73
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__528__B2
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_98
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__528__A2
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__528__A1
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use scs8hd_dfrtp_4  _661_
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_30_143
timestamp 1586364061
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__558__B
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__393__A
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__669__CLK
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _552_
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  FILLER_30_170
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__591__A
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__593__A1N
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_179
timestamp 1586364061
transform 1 0 17572 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__593__A2N
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_183
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__679__RESETB
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__679__CLK
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_194
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_1  _371_
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__588__A
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__609__B
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__684__CLK
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_dfrtp_4  _684_
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_30_252
timestamp 1586364061
transform 1 0 24288 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_240
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 24656 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_xor2_4  _487_
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_31_37
timestamp 1586364061
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__487__B
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__B1
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use scs8hd_o22a_4  _499_
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__653__D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_inv_8  _495_
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__653__CLK
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__390__A
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__528__B1
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _390_
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__558__A
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__524__A
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_o22a_4  _528_
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_xor2_4  _558_
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_31_164
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_155
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__384__A
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__590__B
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _384_
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__590__A
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__679__D
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_dfrtp_4  _679_
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 2154 592
use scs8hd_buf_1  _591_
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 590 592
use scs8hd_decap_6  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__596__A
timestamp 1586364061
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__368__A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__A
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _369_
timestamp 1586364061
transform 1 0 21896 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_243
timestamp 1586364061
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 24656 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__A1N
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__649__RESETB
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_8  _481_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__486__B2
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _496_
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_32_52
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__653__RESETB
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use scs8hd_dfrtp_4  _653_
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_90
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__525__A
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _525_
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_8  _524_
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_120
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__670__RESETB
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_1  _393_
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__383__A
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_and2_4  _590_
timestamp 1586364061
transform 1 0 15456 0 -1 20128
box -38 -48 682 592
use scs8hd_decap_4  FILLER_32_189
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__593__B1
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_a2bb2o_4  _593_
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 1510 592
use scs8hd_decap_8  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_195
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__589__A
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_8  _588_
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_232
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_220
timestamp 1586364061
transform 1 0 21344 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__681__CLK
timestamp 1586364061
transform 1 0 21528 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _596_
timestamp 1586364061
transform 1 0 22540 0 -1 20128
box -38 -48 866 592
use scs8hd_buf_1  _368_
timestamp 1586364061
transform 1 0 21068 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_250
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_242
timestamp 1586364061
transform 1 0 23368 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 24656 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_9
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__649__D
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__486__B1
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_dfrtp_4  _649_
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 2154 592
use scs8hd_a2bb2o_4  _486_
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_25
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__649__CLK
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_1  _407_
timestamp 1586364061
transform 1 0 4232 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_37
timestamp 1586364061
transform 1 0 4508 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_42
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_38
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__499__B2
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__407__A
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__654__D
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_dfrtp_4  _654_
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__654__RESETB
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__654__CLK
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_67
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__664__CLK
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__664__D
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_79
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_75
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__663__CLK
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__664__RESETB
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_90
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_86
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__536__B1
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__536__A1N
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfrtp_4  _664_
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 2154 592
use scs8hd_decap_8  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__531__A
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _531_
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 866 592
use scs8hd_buf_1  _391_
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__A
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_118
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__532__A
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  _389_
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__389__A
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__666__RESETB
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__387__A
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _387_
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_133
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__670__D
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _383_
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 314 592
use scs8hd_dfrtp_4  _670_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 2154 592
use scs8hd_decap_8  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_149
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_163
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__670__CLK
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__594__A
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_xor2_4  _594_
timestamp 1586364061
transform 1 0 16008 0 -1 21216
box -38 -48 2062 592
use scs8hd_decap_8  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_167
timestamp 1586364061
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__593__B2
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__594__B
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_184
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__592__B2
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__592__A1
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__592__B1
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_192
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__682__RESETB
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__682__D
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _589_
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__682__CLK
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__601__A
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_dfrtp_4  _682_
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_34_220
timestamp 1586364061
transform 1 0 21344 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_228
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__599__A2
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__681__RESETB
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__681__D
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use scs8hd_dfrtp_4  _681_
timestamp 1586364061
transform 1 0 21528 0 -1 21216
box -38 -48 2154 592
use scs8hd_decap_8  FILLER_34_245
timestamp 1586364061
transform 1 0 23644 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 24656 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 24656 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__B1
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_o22a_4  _485_
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__485__A2
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _404_
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_42
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__B
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__501__A
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__A
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_46
timestamp 1586364061
transform 1 0 5336 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_58
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_84
timestamp 1586364061
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_80
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__536__B2
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__663__RESETB
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__663__D
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_dfrtp_4  _663_
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 2154 592
use scs8hd_fill_1  FILLER_35_117
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__666__D
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_dfrtp_4  _666_
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_35_165
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_152
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__546__A
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__A
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__386__A
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__680__RESETB
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_181
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__680__D
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_o22a_4  _592_
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_35_213
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_209
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_200
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__592__A2
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__370__A
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _370_
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_217
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__599__A1
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__599__B1
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use scs8hd_o22a_4  _599_
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 1326 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 24656 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_11
timestamp 1586364061
transform 1 0 2116 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__484__A
timestamp 1586364061
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__A1
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_8  _482_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__482__A
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__485__B2
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_xor2_4  _501_
timestamp 1586364061
transform 1 0 4692 0 -1 22304
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_36_71
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_61
timestamp 1586364061
transform 1 0 6716 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__537__A
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_6  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__537__B
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__477__A
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_90
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__536__A2N
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_a2bb2o_4  _536_
timestamp 1586364061
transform 1 0 9844 0 -1 22304
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_36_115
timestamp 1586364061
transform 1 0 11684 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__A2
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _532_
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_130
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_126
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__666__CLK
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__668__CLK
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__668__RESETB
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _385_
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_159
timestamp 1586364061
transform 1 0 15732 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__B2
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__667__CLK
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__667__RESETB
timestamp 1586364061
transform 1 0 15916 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_180
timestamp 1586364061
transform 1 0 17664 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_177
timestamp 1586364061
transform 1 0 17388 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_171
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__680__CLK
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use scs8hd_dfrtp_4  _680_
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 2154 592
use scs8hd_buf_1  _386_
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_212
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_209
timestamp 1586364061
transform 1 0 20332 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_205
timestamp 1586364061
transform 1 0 19964 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__601__B
timestamp 1586364061
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use scs8hd_xor2_4  _601_
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_243
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__599__B2
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 24656 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_9
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__652__D
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_dfrtp_4  _652_
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 2154 592
use scs8hd_decap_3  FILLER_37_45
timestamp 1586364061
transform 1 0 5244 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_41
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_38
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__651__RESETB
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__651__D
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__651__CLK
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__405__A
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _405_
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_67
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__498__A
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_xor2_4  _537_
timestamp 1586364061
transform 1 0 7452 0 1 22304
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_37_91
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__535__B1
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__B1
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_o22a_4  _535_
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__668__D
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_dfrtp_4  _668_
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_155
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__667__D
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _546_
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_181
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_177
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__677__CLK
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__677__RESETB
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_dfrtp_4  _677_
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_37_211
timestamp 1586364061
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_218
timestamp 1586364061
transform 1 0 21160 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_215
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__600__A1N
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__595__A
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_a2bb2o_4  _600_
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1510 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_decap_4  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 24656 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_8
timestamp 1586364061
transform 1 0 1840 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  _484_
timestamp 1586364061
transform 1 0 1564 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_17
timestamp 1586364061
transform 1 0 2668 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_13
timestamp 1586364061
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__494__A
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__652__RESETB
timestamp 1586364061
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_21
timestamp 1586364061
transform 1 0 3036 0 -1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__652__CLK
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_37
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__B2
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_dfrtp_4  _651_
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 2154 592
use scs8hd_decap_4  FILLER_38_66
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_62
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__A1
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _498_
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_90
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_73
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__534__A
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_1  _534_
timestamp 1586364061
transform 1 0 9844 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  _477_
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_98
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__535__A2
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__535__A1
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_116
timestamp 1586364061
transform 1 0 11776 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__535__B2
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__542__A1
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 222 592
use scs8hd_o22a_4  _542_
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_136
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__665__CLK
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__B1
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__A1N
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_151
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_148
timestamp 1586364061
transform 1 0 14720 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__550__A2N
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__A1N
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_dfrtp_4  _667_
timestamp 1586364061
transform 1 0 15916 0 -1 23392
box -38 -48 2154 592
use scs8hd_fill_2  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_184
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__677__D
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_198
timestamp 1586364061
transform 1 0 19320 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_194
timestamp 1586364061
transform 1 0 18952 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__B2
timestamp 1586364061
transform 1 0 19872 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__A2
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__586__A2N
timestamp 1586364061
transform 1 0 18768 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__A1
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_230
timestamp 1586364061
transform 1 0 22264 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_226
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_222
timestamp 1586364061
transform 1 0 21528 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_219
timestamp 1586364061
transform 1 0 21252 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__600__B2
timestamp 1586364061
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__600__B1
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__600__A2N
timestamp 1586364061
transform 1 0 21344 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_8  _595_
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_245
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 24656 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__483__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__483__B
timestamp 1586364061
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_and2_4  _483_
timestamp 1586364061
transform 1 0 1564 0 -1 24480
box -38 -48 682 592
use scs8hd_decap_3  FILLER_40_12
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__494__B
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_17
timestamp 1586364061
transform 1 0 2668 0 -1 24480
box -38 -48 1142 592
use scs8hd_xor2_4  _494_
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 2062 592
use scs8hd_decap_4  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_29
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_41
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_37
timestamp 1586364061
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__B1
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__A2N
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__493__A1N
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use scs8hd_a2bb2o_4  _493_
timestamp 1586364061
transform 1 0 4416 0 -1 24480
box -38 -48 1510 592
use scs8hd_fill_2  FILLER_40_58
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_52
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_49
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__489__A
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__A2
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__B1
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_69
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__492__B2
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_inv_8  _489_
timestamp 1586364061
transform 1 0 6624 0 -1 24480
box -38 -48 866 592
use scs8hd_o22a_4  _492_
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_and2_4  _540_
timestamp 1586364061
transform 1 0 8188 0 -1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__540__A
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__476__A
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__540__B
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_95
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_1  _541_
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_103
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__B
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__544__A
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__541__A
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_112
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__B2
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__543__A2N
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__665__D
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_xor2_4  _544_
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 2062 592
use scs8hd_fill_2  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_120
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__665__RESETB
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_dfrtp_4  _665_
timestamp 1586364061
transform 1 0 12604 0 1 23392
box -38 -48 2154 592
use scs8hd_a2bb2o_4  _543_
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 1510 592
use scs8hd_decap_4  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_147
timestamp 1586364061
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_148
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__549__B2
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__B1
timestamp 1586364061
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__B1
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 130 592
use scs8hd_a2bb2o_4  _550_
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 1510 592
use scs8hd_o22a_4  _549_
timestamp 1586364061
transform 1 0 15732 0 -1 24480
box -38 -48 1326 592
use scs8hd_decap_4  FILLER_40_177
timestamp 1586364061
transform 1 0 17388 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_173
timestamp 1586364061
transform 1 0 17020 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_176
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_172
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__550__B2
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__A2
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__549__A1
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_181
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__586__B2
timestamp 1586364061
transform 1 0 17848 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_184
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__586__B1
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__586__A1N
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_a2bb2o_4  _586_
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1510 592
use scs8hd_decap_8  FILLER_40_206
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_194
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__581__A
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__585__B1
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_o22a_4  _585_
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1326 592
use scs8hd_fill_2  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_inv_8  _582_
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 866 592
use scs8hd_inv_8  _581_
timestamp 1586364061
transform 1 0 21068 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_232
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_226
timestamp 1586364061
transform 1 0 21896 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_231
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__582__A
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__583__B
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_and2_4  _583_
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 682 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__583__A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_252
timestamp 1586364061
transform 1 0 24288 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_240
timestamp 1586364061
transform 1 0 23184 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 24656 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 24656 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_42
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_31
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__491__A
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__490__B
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_buf_1  _491_
timestamp 1586364061
transform 1 0 4140 0 1 24480
box -38 -48 314 592
use scs8hd_inv_8  _488_
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_69
timestamp 1586364061
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_66
timestamp 1586364061
transform 1 0 7176 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__497__A
timestamp 1586364061
transform 1 0 7268 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__488__A
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__497__B
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_82
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_73
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__476__B
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_and2_4  _533_
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 682 592
use scs8hd_and2_4  _497_
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 682 592
use scs8hd_decap_4  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_41_101
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_97
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__547__B
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__533__B
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_inv_8  _538_
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_120
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__547__A
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_xor2_4  _551_
timestamp 1586364061
transform 1 0 13892 0 1 24480
box -38 -48 2062 592
use scs8hd_and2_4  _547_
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 682 592
use scs8hd_decap_4  FILLER_41_165
timestamp 1586364061
transform 1 0 16284 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_161
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__548__A
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_181
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_177
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__587__B
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__587__A
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__545__A
timestamp 1586364061
transform 1 0 16652 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_xor2_4  _587_
timestamp 1586364061
transform 1 0 18216 0 1 24480
box -38 -48 2062 592
use scs8hd_decap_6  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__584__A
timestamp 1586364061
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_227
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_221
timestamp 1586364061
transform 1 0 21436 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_216
timestamp 1586364061
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__597__A
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__597__B
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_and2_4  _597_
timestamp 1586364061
transform 1 0 22172 0 1 24480
box -38 -48 682 592
use scs8hd_buf_1  _584_
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 24656 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_40
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_and2_4  _490_
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 682 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_60
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_52
timestamp 1586364061
transform 1 0 5888 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_48
timestamp 1586364061
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__490__A
timestamp 1586364061
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_and2_4  _476_
timestamp 1586364061
transform 1 0 8280 0 -1 25568
box -38 -48 682 592
use scs8hd_fill_1  FILLER_42_119
timestamp 1586364061
transform 1 0 12052 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_107
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_42_104
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_98
timestamp 1586364061
transform 1 0 10120 0 -1 25568
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__533__A
timestamp 1586364061
transform 1 0 9936 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__538__A
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_142
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_122
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__539__A
timestamp 1586364061
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__551__A
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_8  _539_
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_161
timestamp 1586364061
transform 1 0 15916 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_146
timestamp 1586364061
transform 1 0 14536 0 -1 25568
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__551__B
timestamp 1586364061
transform 1 0 14352 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_1  _548_
timestamp 1586364061
transform 1 0 15640 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_8  _545_
timestamp 1586364061
transform 1 0 16652 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_238
timestamp 1586364061
transform 1 0 23000 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_234
timestamp 1586364061
transform 1 0 22632 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__598__A
timestamp 1586364061
transform 1 0 22816 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_buf_1  _598_
timestamp 1586364061
transform 1 0 22356 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_246
timestamp 1586364061
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 24656 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 20810 27171 20866 27971 6 clk
port 0 nsew default input
rlabel metal2 s 14830 0 14886 800 6 p
port 1 nsew default tristate
rlabel metal2 s 2410 0 2466 800 6 rst
port 2 nsew default input
rlabel metal2 s 18 0 74 800 6 x[0]
port 3 nsew default input
rlabel metal3 s 0 7216 800 7336 6 x[10]
port 4 nsew default input
rlabel metal2 s 22282 0 22338 800 6 x[11]
port 5 nsew default input
rlabel metal3 s 25027 2184 25827 2304 6 x[12]
port 6 nsew default input
rlabel metal2 s 7378 0 7434 800 6 x[13]
port 7 nsew default input
rlabel metal2 s 10874 27171 10930 27971 6 x[14]
port 8 nsew default input
rlabel metal2 s 3422 27171 3478 27971 6 x[15]
port 9 nsew default input
rlabel metal2 s 15842 27171 15898 27971 6 x[16]
port 10 nsew default input
rlabel metal3 s 0 14560 800 14680 6 x[17]
port 11 nsew default input
rlabel metal3 s 25027 5856 25827 5976 6 x[18]
port 12 nsew default input
rlabel metal2 s 24766 0 24822 800 6 x[19]
port 13 nsew default input
rlabel metal3 s 0 10888 800 11008 6 x[1]
port 14 nsew default input
rlabel metal2 s 4894 0 4950 800 6 x[20]
port 15 nsew default input
rlabel metal3 s 25027 24216 25827 24336 6 x[21]
port 16 nsew default input
rlabel metal3 s 0 18232 800 18352 6 x[22]
port 17 nsew default input
rlabel metal2 s 23294 27171 23350 27971 6 x[23]
port 18 nsew default input
rlabel metal2 s 8390 27171 8446 27971 6 x[24]
port 19 nsew default input
rlabel metal3 s 25027 20544 25827 20664 6 x[25]
port 20 nsew default input
rlabel metal2 s 19798 0 19854 800 6 x[26]
port 21 nsew default input
rlabel metal3 s 0 21904 800 22024 6 x[27]
port 22 nsew default input
rlabel metal3 s 25027 16872 25827 16992 6 x[28]
port 23 nsew default input
rlabel metal3 s 0 3544 800 3664 6 x[29]
port 24 nsew default input
rlabel metal2 s 12346 0 12402 800 6 x[2]
port 25 nsew default input
rlabel metal3 s 25027 9528 25827 9648 6 x[30]
port 26 nsew default input
rlabel metal3 s 25027 13200 25827 13320 6 x[31]
port 27 nsew default input
rlabel metal2 s 938 27171 994 27971 6 x[3]
port 28 nsew default input
rlabel metal2 s 18326 27171 18382 27971 6 x[4]
port 29 nsew default input
rlabel metal2 s 17314 0 17370 800 6 x[5]
port 30 nsew default input
rlabel metal2 s 13358 27171 13414 27971 6 x[6]
port 31 nsew default input
rlabel metal3 s 0 25576 800 25696 6 x[7]
port 32 nsew default input
rlabel metal2 s 5906 27171 5962 27971 6 x[8]
port 33 nsew default input
rlabel metal2 s 25686 27171 25742 27971 6 x[9]
port 34 nsew default input
rlabel metal2 s 9862 0 9918 800 6 y
port 35 nsew default input
rlabel metal5 s 1104 5298 24656 5618 6 VDD
port 36 nsew default input
rlabel metal5 s 1104 20616 24656 20936 6 VSS
port 37 nsew default input
<< properties >>
string FIXED_BBOX 0 0 25827 27971
<< end >>
