module spm (clk,
    p,
    rst,
    y,
    VDD,
    VSS,
    x);
 input clk;
 output p;
 input rst;
 input y;
 input VDD;
 input VSS;
 input [31:0] x;

 scs8hd_and2_4 _331_ (.A(_297_),
    .B(x[28]),
    .X(_318_));
 scs8hd_buf_1 _332_ (.A(_318_),
    .X(_319_));
 scs8hd_o22a_4 _333_ (.A2(_317_),
    .A1(_316_),
    .X(_320_),
    .B1(_082_),
    .B2(\pp[29] ));
 scs8hd_a2bb2o_4 _334_ (.A2N(_317_),
    .A1N(_316_),
    .X(_038_),
    .B2(_320_),
    .B1(_319_));
 scs8hd_xor2_4 _335_ (.A(_319_),
    .B(_320_),
    .X(_039_));
 scs8hd_inv_8 _336_ (.Y(_321_),
    .A(_083_));
 scs8hd_inv_8 _337_ (.Y(_322_),
    .A(\pp[30] ));
 scs8hd_and2_4 _338_ (.A(_297_),
    .B(x[29]),
    .X(_323_));
 scs8hd_buf_1 _339_ (.A(_323_),
    .X(_324_));
 scs8hd_o22a_4 _340_ (.A2(_322_),
    .A1(_321_),
    .X(_325_),
    .B1(_083_),
    .B2(\pp[30] ));
 scs8hd_a2bb2o_4 _341_ (.A2N(_322_),
    .A1N(_321_),
    .X(_040_),
    .B2(_325_),
    .B1(_324_));
 scs8hd_xor2_4 _342_ (.A(_324_),
    .B(_325_),
    .X(_041_));
 scs8hd_inv_8 _343_ (.Y(_326_),
    .A(_085_));
 scs8hd_inv_8 _344_ (.Y(_327_),
    .A(\tcmp.s ));
 scs8hd_and2_4 _345_ (.A(_171_),
    .B(x[30]),
    .X(_328_));
 scs8hd_buf_1 _346_ (.A(_328_),
    .X(_329_));
 scs8hd_o22a_4 _347_ (.A2(_327_),
    .A1(_326_),
    .X(_330_),
    .B1(_085_),
    .B2(\tcmp.s ));
 scs8hd_a2bb2o_4 _348_ (.A2N(_327_),
    .A1N(_326_),
    .X(_044_),
    .B2(_330_),
    .B1(_329_));
 scs8hd_xor2_4 _349_ (.A(_329_),
    .B(_330_),
    .X(_045_));
 scs8hd_buf_1 _350_ (.A(_158_),
    .X(_156_));
 scs8hd_inv_8 _351_ (.Y(_157_),
    .A(rst));
 scs8hd_buf_1 _352_ (.A(_157_),
    .X(_155_));
 scs8hd_buf_1 _353_ (.A(_155_),
    .X(_154_));
 scs8hd_buf_1 _354_ (.A(_155_),
    .X(_153_));
 scs8hd_buf_1 _355_ (.A(_155_),
    .X(_152_));
 scs8hd_buf_1 _356_ (.A(_155_),
    .X(_151_));
 scs8hd_buf_1 _357_ (.A(_155_),
    .X(_150_));
 scs8hd_buf_1 _358_ (.A(_157_),
    .X(_158_));
 scs8hd_buf_1 _359_ (.A(_158_),
    .X(_159_));
 scs8hd_buf_1 _360_ (.A(_159_),
    .X(_149_));
 scs8hd_buf_1 _361_ (.A(_159_),
    .X(_148_));
 scs8hd_buf_1 _362_ (.A(_159_),
    .X(_147_));
 scs8hd_buf_1 _363_ (.A(_159_),
    .X(_146_));
 scs8hd_buf_1 _364_ (.A(_159_),
    .X(_145_));
 scs8hd_buf_1 _365_ (.A(_159_),
    .X(_144_));
 scs8hd_buf_1 _366_ (.A(_158_),
    .X(_160_));
 scs8hd_buf_1 _367_ (.A(_160_),
    .X(_143_));
 scs8hd_buf_1 _368_ (.A(_160_),
    .X(_142_));
 scs8hd_buf_1 _369_ (.A(_160_),
    .X(_141_));
 scs8hd_buf_1 _370_ (.A(_160_),
    .X(_140_));
 scs8hd_buf_1 _371_ (.A(_160_),
    .X(_139_));
 scs8hd_buf_1 _372_ (.A(_160_),
    .X(_138_));
 scs8hd_buf_1 _373_ (.A(_157_),
    .X(_161_));
 scs8hd_buf_1 _374_ (.A(_161_),
    .X(_162_));
 scs8hd_buf_1 _375_ (.A(_162_),
    .X(_137_));
 scs8hd_buf_1 _376_ (.A(_162_),
    .X(_136_));
 scs8hd_buf_1 _377_ (.A(_162_),
    .X(_135_));
 scs8hd_buf_1 _378_ (.A(_162_),
    .X(_134_));
 scs8hd_buf_1 _379_ (.A(_162_),
    .X(_133_));
 scs8hd_buf_1 _380_ (.A(_162_),
    .X(_132_));
 scs8hd_buf_1 _381_ (.A(_161_),
    .X(_163_));
 scs8hd_buf_1 _382_ (.A(_163_),
    .X(_131_));
 scs8hd_buf_1 _383_ (.A(_163_),
    .X(_130_));
 scs8hd_buf_1 _384_ (.A(_163_),
    .X(_129_));
 scs8hd_buf_1 _385_ (.A(_163_),
    .X(_128_));
 scs8hd_buf_1 _386_ (.A(_163_),
    .X(_127_));
 scs8hd_buf_1 _387_ (.A(_163_),
    .X(_126_));
 scs8hd_buf_1 _388_ (.A(_161_),
    .X(_164_));
 scs8hd_buf_1 _389_ (.A(_164_),
    .X(_125_));
 scs8hd_buf_1 _390_ (.A(_164_),
    .X(_124_));
 scs8hd_buf_1 _391_ (.A(_164_),
    .X(_123_));
 scs8hd_buf_1 _392_ (.A(_164_),
    .X(_122_));
 scs8hd_buf_1 _393_ (.A(_164_),
    .X(_121_));
 scs8hd_buf_1 _394_ (.A(_164_),
    .X(_120_));
 scs8hd_buf_1 _395_ (.A(_161_),
    .X(_165_));
 scs8hd_buf_1 _396_ (.A(_165_),
    .X(_119_));
 scs8hd_buf_1 _397_ (.A(_165_),
    .X(_118_));
 scs8hd_buf_1 _398_ (.A(_165_),
    .X(_117_));
 scs8hd_buf_1 _399_ (.A(_165_),
    .X(_116_));
 scs8hd_buf_1 _400_ (.A(_165_),
    .X(_115_));
 scs8hd_buf_1 _401_ (.A(_165_),
    .X(_114_));
 scs8hd_buf_1 _402_ (.A(_161_),
    .X(_166_));
 scs8hd_buf_1 _403_ (.A(_166_),
    .X(_113_));
 scs8hd_buf_1 _404_ (.A(_166_),
    .X(_112_));
 scs8hd_buf_1 _405_ (.A(_166_),
    .X(_111_));
 scs8hd_buf_1 _406_ (.A(_166_),
    .X(_110_));
 scs8hd_buf_1 _407_ (.A(_166_),
    .X(_109_));
 scs8hd_buf_1 _408_ (.A(_166_),
    .X(_108_));
 scs8hd_buf_1 _409_ (.A(_161_),
    .X(_167_));
 scs8hd_buf_1 _410_ (.A(_167_),
    .X(_107_));
 scs8hd_buf_1 _411_ (.A(_167_),
    .X(_106_));
 scs8hd_buf_1 _412_ (.A(_167_),
    .X(_105_));
 scs8hd_buf_1 _413_ (.A(_167_),
    .X(_104_));
 scs8hd_buf_1 _414_ (.A(_167_),
    .X(_103_));
 scs8hd_buf_1 _415_ (.A(_167_),
    .X(_102_));
 scs8hd_buf_1 _416_ (.A(_157_),
    .X(_168_));
 scs8hd_buf_1 _417_ (.A(_168_),
    .X(_101_));
 scs8hd_buf_1 _418_ (.A(_168_),
    .X(_100_));
 scs8hd_buf_1 _419_ (.A(_168_),
    .X(_099_));
 scs8hd_buf_1 _420_ (.A(_168_),
    .X(_098_));
 scs8hd_buf_1 _421_ (.A(_168_),
    .X(_097_));
 scs8hd_buf_1 _422_ (.A(_168_),
    .X(_096_));
 scs8hd_buf_1 _423_ (.A(_158_),
    .X(_095_));
 scs8hd_buf_1 _424_ (.A(_158_),
    .X(_094_));
 scs8hd_buf_1 _425_ (.A(_158_),
    .X(_093_));
 scs8hd_inv_8 _426_ (.Y(_169_),
    .A(\csa0.sc ));
 scs8hd_inv_8 _427_ (.Y(_170_),
    .A(\csa0.y ));
 scs8hd_buf_1 _428_ (.A(y),
    .X(_171_));
 scs8hd_buf_1 _429_ (.A(_171_),
    .X(_172_));
 scs8hd_and2_4 _430_ (.A(_172_),
    .B(x[0]),
    .X(_173_));
 scs8hd_buf_1 _431_ (.A(_173_),
    .X(_174_));
 scs8hd_o22a_4 _432_ (.A2(_170_),
    .A1(_169_),
    .X(_175_),
    .B1(\csa0.sc ),
    .B2(\csa0.y ));
 scs8hd_a2bb2o_4 _433_ (.A2N(_170_),
    .A1N(_169_),
    .X(_060_),
    .B2(_175_),
    .B1(_174_));
 scs8hd_xor2_4 _434_ (.A(_174_),
    .B(_175_),
    .X(\csa0.hsum2 ));
 scs8hd_and2_4 _435_ (.A(_171_),
    .B(x[31]),
    .X(_176_));
 scs8hd_or2_4 _436_ (.B(_176_),
    .A(\tcmp.z ),
    .X(_062_));
 scs8hd_a21boi_4 _437_ (.A2(_176_),
    .B1N(_062_),
    .A1(\tcmp.z ),
    .Y(_061_));
 scs8hd_inv_8 _438_ (.Y(_177_),
    .A(_073_));
 scs8hd_inv_8 _439_ (.Y(_178_),
    .A(\pp[2] ));
 scs8hd_and2_4 _440_ (.A(_172_),
    .B(x[1]),
    .X(_179_));
 scs8hd_buf_1 _441_ (.A(_179_),
    .X(_180_));
 scs8hd_o22a_4 _442_ (.A2(_178_),
    .A1(_177_),
    .X(_181_),
    .B1(_073_),
    .B2(\pp[2] ));
 scs8hd_a2bb2o_4 _443_ (.A2N(_178_),
    .A1N(_177_),
    .X(_020_),
    .B2(_181_),
    .B1(_180_));
 scs8hd_xor2_4 _444_ (.A(_180_),
    .B(_181_),
    .X(_021_));
 scs8hd_inv_8 _445_ (.Y(_182_),
    .A(_084_));
 scs8hd_inv_8 _446_ (.Y(_183_),
    .A(\pp[3] ));
 scs8hd_and2_4 _447_ (.A(_172_),
    .B(x[2]),
    .X(_184_));
 scs8hd_buf_1 _448_ (.A(_184_),
    .X(_185_));
 scs8hd_o22a_4 _449_ (.A2(_183_),
    .A1(_182_),
    .X(_186_),
    .B1(_084_),
    .B2(\pp[3] ));
 scs8hd_a2bb2o_4 _450_ (.A2N(_183_),
    .A1N(_182_),
    .X(_042_),
    .B2(_186_),
    .B1(_185_));
 scs8hd_xor2_4 _451_ (.A(_185_),
    .B(_186_),
    .X(_043_));
 scs8hd_inv_8 _452_ (.Y(_187_),
    .A(_086_));
 scs8hd_inv_8 _453_ (.Y(_188_),
    .A(\pp[4] ));
 scs8hd_and2_4 _454_ (.A(_172_),
    .B(x[3]),
    .X(_189_));
 scs8hd_buf_1 _455_ (.A(_189_),
    .X(_190_));
 scs8hd_o22a_4 _456_ (.A2(_188_),
    .A1(_187_),
    .X(_191_),
    .B1(_086_),
    .B2(\pp[4] ));
 scs8hd_a2bb2o_4 _457_ (.A2N(_188_),
    .A1N(_187_),
    .X(_046_),
    .B2(_191_),
    .B1(_190_));
 scs8hd_xor2_4 _458_ (.A(_190_),
    .B(_191_),
    .X(_047_));
 scs8hd_inv_8 _459_ (.Y(_192_),
    .A(_087_));
 scs8hd_inv_8 _460_ (.Y(_193_),
    .A(\pp[5] ));
 scs8hd_and2_4 _461_ (.A(_172_),
    .B(x[4]),
    .X(_194_));
 scs8hd_buf_1 _462_ (.A(_194_),
    .X(_195_));
 scs8hd_o22a_4 _463_ (.A2(_193_),
    .A1(_192_),
    .X(_196_),
    .B1(_087_),
    .B2(\pp[5] ));
 scs8hd_a2bb2o_4 _464_ (.A2N(_193_),
    .A1N(_192_),
    .X(_048_),
    .B2(_196_),
    .B1(_195_));
 scs8hd_xor2_4 _465_ (.A(_195_),
    .B(_196_),
    .X(_049_));
 scs8hd_inv_8 _466_ (.Y(_197_),
    .A(_088_));
 scs8hd_inv_8 _467_ (.Y(_198_),
    .A(\pp[6] ));
 scs8hd_and2_4 _468_ (.A(_172_),
    .B(x[5]),
    .X(_199_));
 scs8hd_buf_1 _469_ (.A(_199_),
    .X(_200_));
 scs8hd_o22a_4 _470_ (.A2(_198_),
    .A1(_197_),
    .X(_201_),
    .B1(_088_),
    .B2(\pp[6] ));
 scs8hd_a2bb2o_4 _471_ (.A2N(_198_),
    .A1N(_197_),
    .X(_050_),
    .B2(_201_),
    .B1(_200_));
 scs8hd_xor2_4 _472_ (.A(_200_),
    .B(_201_),
    .X(_051_));
 scs8hd_inv_8 _473_ (.Y(_202_),
    .A(_089_));
 scs8hd_inv_8 _474_ (.Y(_203_),
    .A(\pp[7] ));
 scs8hd_buf_1 _475_ (.A(_171_),
    .X(_204_));
 scs8hd_and2_4 _476_ (.A(_204_),
    .B(x[6]),
    .X(_205_));
 scs8hd_buf_1 _477_ (.A(_205_),
    .X(_206_));
 scs8hd_o22a_4 _478_ (.A2(_203_),
    .A1(_202_),
    .X(_207_),
    .B1(_089_),
    .B2(\pp[7] ));
 scs8hd_a2bb2o_4 _479_ (.A2N(_203_),
    .A1N(_202_),
    .X(_052_),
    .B2(_207_),
    .B1(_206_));
 scs8hd_xor2_4 _480_ (.A(_206_),
    .B(_207_),
    .X(_053_));
 scs8hd_inv_8 _481_ (.Y(_208_),
    .A(_090_));
 scs8hd_inv_8 _482_ (.Y(_209_),
    .A(\pp[8] ));
 scs8hd_and2_4 _483_ (.A(_204_),
    .B(x[7]),
    .X(_210_));
 scs8hd_buf_1 _484_ (.A(_210_),
    .X(_211_));
 scs8hd_o22a_4 _485_ (.A2(_209_),
    .A1(_208_),
    .X(_212_),
    .B1(_090_),
    .B2(\pp[8] ));
 scs8hd_a2bb2o_4 _486_ (.A2N(_209_),
    .A1N(_208_),
    .X(_054_),
    .B2(_212_),
    .B1(_211_));
 scs8hd_xor2_4 _487_ (.A(_211_),
    .B(_212_),
    .X(_055_));
 scs8hd_inv_8 _488_ (.Y(_213_),
    .A(_091_));
 scs8hd_inv_8 _489_ (.Y(_214_),
    .A(\pp[9] ));
 scs8hd_and2_4 _490_ (.A(_204_),
    .B(x[8]),
    .X(_215_));
 scs8hd_buf_1 _491_ (.A(_215_),
    .X(_216_));
 scs8hd_o22a_4 _492_ (.A2(_214_),
    .A1(_213_),
    .X(_217_),
    .B1(_091_),
    .B2(\pp[9] ));
 scs8hd_a2bb2o_4 _493_ (.A2N(_214_),
    .A1N(_213_),
    .X(_056_),
    .B2(_217_),
    .B1(_216_));
 scs8hd_xor2_4 _494_ (.A(_216_),
    .B(_217_),
    .X(_057_));
 scs8hd_inv_8 _495_ (.Y(_218_),
    .A(_092_));
 scs8hd_inv_8 _496_ (.Y(_219_),
    .A(\pp[10] ));
 scs8hd_and2_4 _497_ (.A(_204_),
    .B(x[9]),
    .X(_220_));
 scs8hd_buf_1 _498_ (.A(_220_),
    .X(_221_));
 scs8hd_o22a_4 _499_ (.A2(_219_),
    .A1(_218_),
    .X(_222_),
    .B1(_092_),
    .B2(\pp[10] ));
 scs8hd_a2bb2o_4 _500_ (.A2N(_219_),
    .A1N(_218_),
    .X(_058_),
    .B2(_222_),
    .B1(_221_));
 scs8hd_xor2_4 _501_ (.A(_221_),
    .B(_222_),
    .X(_059_));
 scs8hd_inv_8 _502_ (.Y(_223_),
    .A(_063_));
 scs8hd_inv_8 _503_ (.Y(_224_),
    .A(\pp[11] ));
 scs8hd_and2_4 _504_ (.A(_204_),
    .B(x[10]),
    .X(_225_));
 scs8hd_buf_1 _505_ (.A(_225_),
    .X(_226_));
 scs8hd_o22a_4 _506_ (.A2(_224_),
    .A1(_223_),
    .X(_227_),
    .B1(_063_),
    .B2(\pp[11] ));
 scs8hd_a2bb2o_4 _507_ (.A2N(_224_),
    .A1N(_223_),
    .X(_000_),
    .B2(_227_),
    .B1(_226_));
 scs8hd_xor2_4 _508_ (.A(_226_),
    .B(_227_),
    .X(_001_));
 scs8hd_inv_8 _509_ (.Y(_228_),
    .A(_064_));
 scs8hd_inv_8 _510_ (.Y(_229_),
    .A(\pp[12] ));
 scs8hd_and2_4 _511_ (.A(_204_),
    .B(x[11]),
    .X(_230_));
 scs8hd_buf_1 _512_ (.A(_230_),
    .X(_231_));
 scs8hd_o22a_4 _513_ (.A2(_229_),
    .A1(_228_),
    .X(_232_),
    .B1(_064_),
    .B2(\pp[12] ));
 scs8hd_a2bb2o_4 _514_ (.A2N(_229_),
    .A1N(_228_),
    .X(_002_),
    .B2(_232_),
    .B1(_231_));
 scs8hd_xor2_4 _515_ (.A(_231_),
    .B(_232_),
    .X(_003_));
 scs8hd_inv_8 _516_ (.Y(_233_),
    .A(_065_));
 scs8hd_inv_8 _517_ (.Y(_234_),
    .A(\pp[13] ));
 scs8hd_buf_1 _518_ (.A(_171_),
    .X(_235_));
 scs8hd_and2_4 _519_ (.A(_235_),
    .B(x[12]),
    .X(_236_));
 scs8hd_buf_1 _520_ (.A(_236_),
    .X(_237_));
 scs8hd_o22a_4 _521_ (.A2(_234_),
    .A1(_233_),
    .X(_238_),
    .B1(_065_),
    .B2(\pp[13] ));
 scs8hd_a2bb2o_4 _522_ (.A2N(_234_),
    .A1N(_233_),
    .X(_004_),
    .B2(_238_),
    .B1(_237_));
 scs8hd_xor2_4 _523_ (.A(_237_),
    .B(_238_),
    .X(_005_));
 scs8hd_inv_8 _524_ (.Y(_239_),
    .A(_066_));
 scs8hd_inv_8 _525_ (.Y(_240_),
    .A(\pp[14] ));
 scs8hd_and2_4 _526_ (.A(_235_),
    .B(x[13]),
    .X(_241_));
 scs8hd_buf_1 _527_ (.A(_241_),
    .X(_242_));
 scs8hd_o22a_4 _528_ (.A2(_240_),
    .A1(_239_),
    .X(_243_),
    .B1(_066_),
    .B2(\pp[14] ));
 scs8hd_a2bb2o_4 _529_ (.A2N(_240_),
    .A1N(_239_),
    .X(_006_),
    .B2(_243_),
    .B1(_242_));
 scs8hd_xor2_4 _530_ (.A(_242_),
    .B(_243_),
    .X(_007_));
 scs8hd_inv_8 _531_ (.Y(_244_),
    .A(_067_));
 scs8hd_inv_8 _532_ (.Y(_245_),
    .A(\pp[15] ));
 scs8hd_and2_4 _533_ (.A(_235_),
    .B(x[14]),
    .X(_246_));
 scs8hd_buf_1 _534_ (.A(_246_),
    .X(_247_));
 scs8hd_o22a_4 _535_ (.A2(_245_),
    .A1(_244_),
    .X(_248_),
    .B1(_067_),
    .B2(\pp[15] ));
 scs8hd_a2bb2o_4 _536_ (.A2N(_245_),
    .A1N(_244_),
    .X(_008_),
    .B2(_248_),
    .B1(_247_));
 scs8hd_xor2_4 _537_ (.A(_247_),
    .B(_248_),
    .X(_009_));
 scs8hd_inv_8 _538_ (.Y(_249_),
    .A(_068_));
 scs8hd_inv_8 _539_ (.Y(_250_),
    .A(\pp[16] ));
 scs8hd_and2_4 _540_ (.A(_235_),
    .B(x[15]),
    .X(_251_));
 scs8hd_buf_1 _541_ (.A(_251_),
    .X(_252_));
 scs8hd_o22a_4 _542_ (.A2(_250_),
    .A1(_249_),
    .X(_253_),
    .B1(_068_),
    .B2(\pp[16] ));
 scs8hd_a2bb2o_4 _543_ (.A2N(_250_),
    .A1N(_249_),
    .X(_010_),
    .B2(_253_),
    .B1(_252_));
 scs8hd_xor2_4 _544_ (.A(_252_),
    .B(_253_),
    .X(_011_));
 scs8hd_inv_8 _545_ (.Y(_254_),
    .A(_069_));
 scs8hd_inv_8 _546_ (.Y(_255_),
    .A(\pp[17] ));
 scs8hd_and2_4 _547_ (.A(_235_),
    .B(x[16]),
    .X(_256_));
 scs8hd_buf_1 _548_ (.A(_256_),
    .X(_257_));
 scs8hd_o22a_4 _549_ (.A2(_255_),
    .A1(_254_),
    .X(_258_),
    .B1(_069_),
    .B2(\pp[17] ));
 scs8hd_a2bb2o_4 _550_ (.A2N(_255_),
    .A1N(_254_),
    .X(_012_),
    .B2(_258_),
    .B1(_257_));
 scs8hd_xor2_4 _551_ (.A(_257_),
    .B(_258_),
    .X(_013_));
 scs8hd_inv_8 _552_ (.Y(_259_),
    .A(_070_));
 scs8hd_inv_8 _553_ (.Y(_260_),
    .A(\pp[18] ));
 scs8hd_and2_4 _554_ (.A(_235_),
    .B(x[17]),
    .X(_261_));
 scs8hd_buf_1 _555_ (.A(_261_),
    .X(_262_));
 scs8hd_o22a_4 _556_ (.A2(_260_),
    .A1(_259_),
    .X(_263_),
    .B1(_070_),
    .B2(\pp[18] ));
 scs8hd_a2bb2o_4 _557_ (.A2N(_260_),
    .A1N(_259_),
    .X(_014_),
    .B2(_263_),
    .B1(_262_));
 scs8hd_xor2_4 _558_ (.A(_262_),
    .B(_263_),
    .X(_015_));
 scs8hd_inv_8 _559_ (.Y(_264_),
    .A(_071_));
 scs8hd_inv_8 _560_ (.Y(_265_),
    .A(\pp[19] ));
 scs8hd_buf_1 _561_ (.A(_171_),
    .X(_266_));
 scs8hd_and2_4 _562_ (.A(_266_),
    .B(x[18]),
    .X(_267_));
 scs8hd_buf_1 _563_ (.A(_267_),
    .X(_268_));
 scs8hd_o22a_4 _564_ (.A2(_265_),
    .A1(_264_),
    .X(_269_),
    .B1(_071_),
    .B2(\pp[19] ));
 scs8hd_a2bb2o_4 _565_ (.A2N(_265_),
    .A1N(_264_),
    .X(_016_),
    .B2(_269_),
    .B1(_268_));
 scs8hd_xor2_4 _566_ (.A(_268_),
    .B(_269_),
    .X(_017_));
 scs8hd_inv_8 _567_ (.Y(_270_),
    .A(_072_));
 scs8hd_inv_8 _568_ (.Y(_271_),
    .A(\pp[20] ));
 scs8hd_and2_4 _569_ (.A(_266_),
    .B(x[19]),
    .X(_272_));
 scs8hd_buf_1 _570_ (.A(_272_),
    .X(_273_));
 scs8hd_o22a_4 _571_ (.A2(_271_),
    .A1(_270_),
    .X(_274_),
    .B1(_072_),
    .B2(\pp[20] ));
 scs8hd_a2bb2o_4 _572_ (.A2N(_271_),
    .A1N(_270_),
    .X(_018_),
    .B2(_274_),
    .B1(_273_));
 scs8hd_xor2_4 _573_ (.A(_273_),
    .B(_274_),
    .X(_019_));
 scs8hd_inv_8 _574_ (.Y(_275_),
    .A(_074_));
 scs8hd_inv_8 _575_ (.Y(_276_),
    .A(\pp[21] ));
 scs8hd_and2_4 _576_ (.A(_266_),
    .B(x[20]),
    .X(_277_));
 scs8hd_buf_1 _577_ (.A(_277_),
    .X(_278_));
 scs8hd_o22a_4 _578_ (.A2(_276_),
    .A1(_275_),
    .X(_279_),
    .B1(_074_),
    .B2(\pp[21] ));
 scs8hd_a2bb2o_4 _579_ (.A2N(_276_),
    .A1N(_275_),
    .X(_022_),
    .B2(_279_),
    .B1(_278_));
 scs8hd_xor2_4 _580_ (.A(_278_),
    .B(_279_),
    .X(_023_));
 scs8hd_inv_8 _581_ (.Y(_280_),
    .A(_075_));
 scs8hd_inv_8 _582_ (.Y(_281_),
    .A(\pp[22] ));
 scs8hd_and2_4 _583_ (.A(_266_),
    .B(x[21]),
    .X(_282_));
 scs8hd_buf_1 _584_ (.A(_282_),
    .X(_283_));
 scs8hd_o22a_4 _585_ (.A2(_281_),
    .A1(_280_),
    .X(_284_),
    .B1(_075_),
    .B2(\pp[22] ));
 scs8hd_a2bb2o_4 _586_ (.A2N(_281_),
    .A1N(_280_),
    .X(_024_),
    .B2(_284_),
    .B1(_283_));
 scs8hd_xor2_4 _587_ (.A(_283_),
    .B(_284_),
    .X(_025_));
 scs8hd_inv_8 _588_ (.Y(_285_),
    .A(_076_));
 scs8hd_inv_8 _589_ (.Y(_286_),
    .A(\pp[23] ));
 scs8hd_and2_4 _590_ (.A(_266_),
    .B(x[22]),
    .X(_287_));
 scs8hd_buf_1 _591_ (.A(_287_),
    .X(_288_));
 scs8hd_o22a_4 _592_ (.A2(_286_),
    .A1(_285_),
    .X(_289_),
    .B1(_076_),
    .B2(\pp[23] ));
 scs8hd_a2bb2o_4 _593_ (.A2N(_286_),
    .A1N(_285_),
    .X(_026_),
    .B2(_289_),
    .B1(_288_));
 scs8hd_xor2_4 _594_ (.A(_288_),
    .B(_289_),
    .X(_027_));
 scs8hd_inv_8 _595_ (.Y(_290_),
    .A(_077_));
 scs8hd_inv_8 _596_ (.Y(_291_),
    .A(\pp[24] ));
 scs8hd_and2_4 _597_ (.A(_266_),
    .B(x[23]),
    .X(_292_));
 scs8hd_buf_1 _598_ (.A(_292_),
    .X(_293_));
 scs8hd_o22a_4 _599_ (.A2(_291_),
    .A1(_290_),
    .X(_294_),
    .B1(_077_),
    .B2(\pp[24] ));
 scs8hd_a2bb2o_4 _600_ (.A2N(_291_),
    .A1N(_290_),
    .X(_028_),
    .B2(_294_),
    .B1(_293_));
 scs8hd_xor2_4 _601_ (.A(_293_),
    .B(_294_),
    .X(_029_));
 scs8hd_inv_8 _602_ (.Y(_295_),
    .A(_078_));
 scs8hd_inv_8 _603_ (.Y(_296_),
    .A(\pp[25] ));
 scs8hd_buf_1 _604_ (.A(y),
    .X(_297_));
 scs8hd_and2_4 _605_ (.A(_297_),
    .B(x[24]),
    .X(_298_));
 scs8hd_buf_1 _606_ (.A(_298_),
    .X(_299_));
 scs8hd_o22a_4 _607_ (.A2(_296_),
    .A1(_295_),
    .X(_300_),
    .B1(_078_),
    .B2(\pp[25] ));
 scs8hd_a2bb2o_4 _608_ (.A2N(_296_),
    .A1N(_295_),
    .X(_030_),
    .B2(_300_),
    .B1(_299_));
 scs8hd_xor2_4 _609_ (.A(_299_),
    .B(_300_),
    .X(_031_));
 scs8hd_inv_8 _610_ (.Y(_301_),
    .A(_079_));
 scs8hd_inv_8 _611_ (.Y(_302_),
    .A(\pp[26] ));
 scs8hd_and2_4 _612_ (.A(_297_),
    .B(x[25]),
    .X(_303_));
 scs8hd_buf_1 _613_ (.A(_303_),
    .X(_304_));
 scs8hd_o22a_4 _614_ (.A2(_302_),
    .A1(_301_),
    .X(_305_),
    .B1(_079_),
    .B2(\pp[26] ));
 scs8hd_a2bb2o_4 _615_ (.A2N(_302_),
    .A1N(_301_),
    .X(_032_),
    .B2(_305_),
    .B1(_304_));
 scs8hd_xor2_4 _616_ (.A(_304_),
    .B(_305_),
    .X(_033_));
 scs8hd_inv_8 _617_ (.Y(_306_),
    .A(_080_));
 scs8hd_inv_8 _618_ (.Y(_307_),
    .A(\pp[27] ));
 scs8hd_and2_4 _619_ (.A(_297_),
    .B(x[26]),
    .X(_308_));
 scs8hd_buf_1 _620_ (.A(_308_),
    .X(_309_));
 scs8hd_o22a_4 _621_ (.A2(_307_),
    .A1(_306_),
    .X(_310_),
    .B1(_080_),
    .B2(\pp[27] ));
 scs8hd_a2bb2o_4 _622_ (.A2N(_307_),
    .A1N(_306_),
    .X(_034_),
    .B2(_310_),
    .B1(_309_));
 scs8hd_xor2_4 _623_ (.A(_309_),
    .B(_310_),
    .X(_035_));
 scs8hd_inv_8 _624_ (.Y(_311_),
    .A(_081_));
 scs8hd_inv_8 _625_ (.Y(_312_),
    .A(\pp[28] ));
 scs8hd_and2_4 _626_ (.A(_297_),
    .B(x[27]),
    .X(_313_));
 scs8hd_buf_1 _627_ (.A(_313_),
    .X(_314_));
 scs8hd_o22a_4 _628_ (.A2(_312_),
    .A1(_311_),
    .X(_315_),
    .B1(_081_),
    .B2(\pp[28] ));
 scs8hd_a2bb2o_4 _629_ (.A2N(_312_),
    .A1N(_311_),
    .X(_036_),
    .B2(_315_),
    .B1(_314_));
 scs8hd_xor2_4 _630_ (.A(_314_),
    .B(_315_),
    .X(_037_));
 scs8hd_inv_8 _631_ (.Y(_316_),
    .A(_082_));
 scs8hd_inv_8 _632_ (.Y(_317_),
    .A(\pp[29] ));
 scs8hd_dfrtp_4 _633_ (.CLK(clk_0_0),
    .D(_060_),
    .RESETB(_093_),
    .Q(\csa0.sc ));
 scs8hd_dfrtp_4 _634_ (.CLK(clk_0_0),
    .D(\csa0.hsum2 ),
    .RESETB(_094_),
    .Q(p));
 scs8hd_dfrtp_4 _635_ (.CLK(clk_0_0),
    .D(_062_),
    .RESETB(_095_),
    .Q(\tcmp.z ));
 scs8hd_dfrtp_4 _636_ (.CLK(clk_0_0),
    .D(_061_),
    .RESETB(_096_),
    .Q(\tcmp.s ));
 scs8hd_dfrtp_4 _637_ (.CLK(clk_0_0),
    .D(_020_),
    .RESETB(_097_),
    .Q(_073_));
 scs8hd_dfrtp_4 _638_ (.CLK(clk_0_0),
    .D(_021_),
    .RESETB(_098_),
    .Q(\csa0.y ));
 scs8hd_dfrtp_4 _639_ (.CLK(clk_0_0),
    .D(_042_),
    .RESETB(_099_),
    .Q(_084_));
 scs8hd_dfrtp_4 _640_ (.CLK(clk_0_0),
    .D(_043_),
    .RESETB(_100_),
    .Q(\pp[2] ));
 scs8hd_dfrtp_4 _641_ (.CLK(clk_0_0),
    .D(_046_),
    .RESETB(_101_),
    .Q(_086_));
 scs8hd_dfrtp_4 _642_ (.CLK(clk_0_0),
    .D(_047_),
    .RESETB(_102_),
    .Q(\pp[3] ));
 scs8hd_dfrtp_4 _643_ (.CLK(clk_0_0),
    .D(_048_),
    .RESETB(_103_),
    .Q(_087_));
 scs8hd_dfrtp_4 _644_ (.CLK(clk_0_0),
    .D(_049_),
    .RESETB(_104_),
    .Q(\pp[4] ));
 scs8hd_dfrtp_4 _645_ (.CLK(clk_0_0),
    .D(_050_),
    .RESETB(_105_),
    .Q(_088_));
 scs8hd_dfrtp_4 _646_ (.CLK(clk_0_0),
    .D(_051_),
    .RESETB(_106_),
    .Q(\pp[5] ));
 scs8hd_dfrtp_4 _647_ (.CLK(clk_0_0),
    .D(_052_),
    .RESETB(_107_),
    .Q(_089_));
 scs8hd_dfrtp_4 _648_ (.CLK(clk_0_0),
    .D(_053_),
    .RESETB(_108_),
    .Q(\pp[6] ));
 scs8hd_dfrtp_4 _649_ (.CLK(clk_0_16),
    .D(_054_),
    .RESETB(_109_),
    .Q(_090_));
 scs8hd_dfrtp_4 _650_ (.CLK(clk_0_16),
    .D(_055_),
    .RESETB(_110_),
    .Q(\pp[7] ));
 scs8hd_dfrtp_4 _651_ (.CLK(clk_0_16),
    .D(_056_),
    .RESETB(_111_),
    .Q(_091_));
 scs8hd_dfrtp_4 _652_ (.CLK(clk_0_16),
    .D(_057_),
    .RESETB(_112_),
    .Q(\pp[8] ));
 scs8hd_dfrtp_4 _653_ (.CLK(clk_0_16),
    .D(_058_),
    .RESETB(_113_),
    .Q(_092_));
 scs8hd_dfrtp_4 _654_ (.CLK(clk_0_16),
    .D(_059_),
    .RESETB(_114_),
    .Q(\pp[9] ));
 scs8hd_dfrtp_4 _655_ (.CLK(clk_0_16),
    .D(_000_),
    .RESETB(_115_),
    .Q(_063_));
 scs8hd_dfrtp_4 _656_ (.CLK(clk_0_16),
    .D(_001_),
    .RESETB(_116_),
    .Q(\pp[10] ));
 scs8hd_dfrtp_4 _657_ (.CLK(clk_0_16),
    .D(_002_),
    .RESETB(_117_),
    .Q(_064_));
 scs8hd_dfrtp_4 _658_ (.CLK(clk_0_16),
    .D(_003_),
    .RESETB(_118_),
    .Q(\pp[11] ));
 scs8hd_dfrtp_4 _659_ (.CLK(clk_0_16),
    .D(_004_),
    .RESETB(_119_),
    .Q(_065_));
 scs8hd_dfrtp_4 _660_ (.CLK(clk_0_16),
    .D(_005_),
    .RESETB(_120_),
    .Q(\pp[12] ));
 scs8hd_dfrtp_4 _661_ (.CLK(clk_0_16),
    .D(_006_),
    .RESETB(_121_),
    .Q(_066_));
 scs8hd_dfrtp_4 _662_ (.CLK(clk_0_16),
    .D(_007_),
    .RESETB(_122_),
    .Q(\pp[13] ));
 scs8hd_dfrtp_4 _663_ (.CLK(clk_0_16),
    .D(_008_),
    .RESETB(_123_),
    .Q(_067_));
 scs8hd_dfrtp_4 _664_ (.CLK(clk_0_16),
    .D(_009_),
    .RESETB(_124_),
    .Q(\pp[14] ));
 scs8hd_dfrtp_4 _665_ (.CLK(clk_0_32),
    .D(_010_),
    .RESETB(_125_),
    .Q(_068_));
 scs8hd_dfrtp_4 _666_ (.CLK(clk_0_32),
    .D(_011_),
    .RESETB(_126_),
    .Q(\pp[15] ));
 scs8hd_dfrtp_4 _667_ (.CLK(clk_0_32),
    .D(_012_),
    .RESETB(_127_),
    .Q(_069_));
 scs8hd_dfrtp_4 _668_ (.CLK(clk_0_32),
    .D(_013_),
    .RESETB(_128_),
    .Q(\pp[16] ));
 scs8hd_dfrtp_4 _669_ (.CLK(clk_0_32),
    .D(_014_),
    .RESETB(_129_),
    .Q(_070_));
 scs8hd_dfrtp_4 _670_ (.CLK(clk_0_32),
    .D(_015_),
    .RESETB(_130_),
    .Q(\pp[17] ));
 scs8hd_dfrtp_4 _671_ (.CLK(clk_0_32),
    .D(_016_),
    .RESETB(_131_),
    .Q(_071_));
 scs8hd_dfrtp_4 _672_ (.CLK(clk_0_32),
    .D(_017_),
    .RESETB(_132_),
    .Q(\pp[18] ));
 scs8hd_dfrtp_4 _673_ (.CLK(clk_0_32),
    .D(_018_),
    .RESETB(_133_),
    .Q(_072_));
 scs8hd_dfrtp_4 _674_ (.CLK(clk_0_32),
    .D(_019_),
    .RESETB(_134_),
    .Q(\pp[19] ));
 scs8hd_dfrtp_4 _675_ (.CLK(clk_0_32),
    .D(_022_),
    .RESETB(_135_),
    .Q(_074_));
 scs8hd_dfrtp_4 _676_ (.CLK(clk_0_32),
    .D(_023_),
    .RESETB(_136_),
    .Q(\pp[20] ));
 scs8hd_dfrtp_4 _677_ (.CLK(clk_0_32),
    .D(_024_),
    .RESETB(_137_),
    .Q(_075_));
 scs8hd_dfrtp_4 _678_ (.CLK(clk_0_32),
    .D(_025_),
    .RESETB(_138_),
    .Q(\pp[21] ));
 scs8hd_dfrtp_4 _679_ (.CLK(clk_0_32),
    .D(_026_),
    .RESETB(_139_),
    .Q(_076_));
 scs8hd_dfrtp_4 _680_ (.CLK(clk_0_32),
    .D(_027_),
    .RESETB(_140_),
    .Q(\pp[22] ));
 scs8hd_dfrtp_4 _681_ (.CLK(clk_0_48),
    .D(_028_),
    .RESETB(_141_),
    .Q(_077_));
 scs8hd_dfrtp_4 _682_ (.CLK(clk_0_48),
    .D(_029_),
    .RESETB(_142_),
    .Q(\pp[23] ));
 scs8hd_dfrtp_4 _683_ (.CLK(clk_0_48),
    .D(_030_),
    .RESETB(_143_),
    .Q(_078_));
 scs8hd_dfrtp_4 _684_ (.CLK(clk_0_48),
    .D(_031_),
    .RESETB(_144_),
    .Q(\pp[24] ));
 scs8hd_dfrtp_4 _685_ (.CLK(clk_0_48),
    .D(_032_),
    .RESETB(_145_),
    .Q(_079_));
 scs8hd_dfrtp_4 _686_ (.CLK(clk_0_48),
    .D(_033_),
    .RESETB(_146_),
    .Q(\pp[25] ));
 scs8hd_dfrtp_4 _687_ (.CLK(clk_0_48),
    .D(_034_),
    .RESETB(_147_),
    .Q(_080_));
 scs8hd_dfrtp_4 _688_ (.CLK(clk_0_48),
    .D(_035_),
    .RESETB(_148_),
    .Q(\pp[26] ));
 scs8hd_dfrtp_4 _689_ (.CLK(clk_0_48),
    .D(_036_),
    .RESETB(_149_),
    .Q(_081_));
 scs8hd_dfrtp_4 _690_ (.CLK(clk_0_48),
    .D(_037_),
    .RESETB(_150_),
    .Q(\pp[27] ));
 scs8hd_dfrtp_4 _691_ (.CLK(clk_0_48),
    .D(_038_),
    .RESETB(_151_),
    .Q(_082_));
 scs8hd_dfrtp_4 _692_ (.CLK(clk_0_48),
    .D(_039_),
    .RESETB(_152_),
    .Q(\pp[28] ));
 scs8hd_dfrtp_4 _693_ (.CLK(clk_0_48),
    .D(_040_),
    .RESETB(_153_),
    .Q(_083_));
 scs8hd_dfrtp_4 _694_ (.CLK(clk_0_48),
    .D(_041_),
    .RESETB(_154_),
    .Q(\pp[29] ));
 scs8hd_dfrtp_4 _695_ (.CLK(clk_0_48),
    .D(_044_),
    .RESETB(_155_),
    .Q(_085_));
 scs8hd_dfrtp_4 _696_ (.CLK(clk_0_48),
    .D(_045_),
    .RESETB(_156_),
    .Q(\pp[30] ));
 scs8hd_clkbuf_4 _CTS_buf_1_0 (.A(clk_1_0),
    .X(clk_0_0));
 scs8hd_clkbuf_4 _CTS_buf_1_16 (.A(clk_1_0),
    .X(clk_0_16));
 scs8hd_clkbuf_4 _CTS_buf_1_32 (.A(clk_1_0),
    .X(clk_0_32));
 scs8hd_clkbuf_4 _CTS_buf_1_48 (.A(clk_1_0),
    .X(clk_0_48));
 scs8hd_clkbuf_16 _CTS_root (.A(clk),
    .X(clk_1_0));
 scs8hd_decap_3 PHY_0 ();
 scs8hd_decap_3 PHY_1 ();
 scs8hd_decap_3 PHY_2 ();
 scs8hd_decap_3 PHY_3 ();
 scs8hd_decap_3 PHY_4 ();
 scs8hd_decap_3 PHY_5 ();
 scs8hd_decap_3 PHY_6 ();
 scs8hd_decap_3 PHY_7 ();
 scs8hd_decap_3 PHY_8 ();
 scs8hd_decap_3 PHY_9 ();
 scs8hd_decap_3 PHY_10 ();
 scs8hd_decap_3 PHY_11 ();
 scs8hd_decap_3 PHY_12 ();
 scs8hd_decap_3 PHY_13 ();
 scs8hd_decap_3 PHY_14 ();
 scs8hd_decap_3 PHY_15 ();
 scs8hd_decap_3 PHY_16 ();
 scs8hd_decap_3 PHY_17 ();
 scs8hd_decap_3 PHY_18 ();
 scs8hd_decap_3 PHY_19 ();
 scs8hd_decap_3 PHY_20 ();
 scs8hd_decap_3 PHY_21 ();
 scs8hd_decap_3 PHY_22 ();
 scs8hd_decap_3 PHY_23 ();
 scs8hd_decap_3 PHY_24 ();
 scs8hd_decap_3 PHY_25 ();
 scs8hd_decap_3 PHY_26 ();
 scs8hd_decap_3 PHY_27 ();
 scs8hd_decap_3 PHY_28 ();
 scs8hd_decap_3 PHY_29 ();
 scs8hd_decap_3 PHY_30 ();
 scs8hd_decap_3 PHY_31 ();
 scs8hd_decap_3 PHY_32 ();
 scs8hd_decap_3 PHY_33 ();
 scs8hd_decap_3 PHY_34 ();
 scs8hd_decap_3 PHY_35 ();
 scs8hd_decap_3 PHY_36 ();
 scs8hd_decap_3 PHY_37 ();
 scs8hd_decap_3 PHY_38 ();
 scs8hd_decap_3 PHY_39 ();
 scs8hd_decap_3 PHY_40 ();
 scs8hd_decap_3 PHY_41 ();
 scs8hd_decap_3 PHY_42 ();
 scs8hd_decap_3 PHY_43 ();
 scs8hd_decap_3 PHY_44 ();
 scs8hd_decap_3 PHY_45 ();
 scs8hd_decap_3 PHY_46 ();
 scs8hd_decap_3 PHY_47 ();
 scs8hd_decap_3 PHY_48 ();
 scs8hd_decap_3 PHY_49 ();
 scs8hd_decap_3 PHY_50 ();
 scs8hd_decap_3 PHY_51 ();
 scs8hd_decap_3 PHY_52 ();
 scs8hd_decap_3 PHY_53 ();
 scs8hd_decap_3 PHY_54 ();
 scs8hd_decap_3 PHY_55 ();
 scs8hd_decap_3 PHY_56 ();
 scs8hd_decap_3 PHY_57 ();
 scs8hd_decap_3 PHY_58 ();
 scs8hd_decap_3 PHY_59 ();
 scs8hd_decap_3 PHY_60 ();
 scs8hd_decap_3 PHY_61 ();
 scs8hd_decap_3 PHY_62 ();
 scs8hd_decap_3 PHY_63 ();
 scs8hd_decap_3 PHY_64 ();
 scs8hd_decap_3 PHY_65 ();
 scs8hd_decap_3 PHY_66 ();
 scs8hd_decap_3 PHY_67 ();
 scs8hd_decap_3 PHY_68 ();
 scs8hd_decap_3 PHY_69 ();
 scs8hd_decap_3 PHY_70 ();
 scs8hd_decap_3 PHY_71 ();
 scs8hd_decap_3 PHY_72 ();
 scs8hd_decap_3 PHY_73 ();
 scs8hd_decap_3 PHY_74 ();
 scs8hd_decap_3 PHY_75 ();
 scs8hd_decap_3 PHY_76 ();
 scs8hd_decap_3 PHY_77 ();
 scs8hd_decap_3 PHY_78 ();
 scs8hd_decap_3 PHY_79 ();
 scs8hd_decap_3 PHY_80 ();
 scs8hd_decap_3 PHY_81 ();
 scs8hd_decap_3 PHY_82 ();
 scs8hd_decap_3 PHY_83 ();
 scs8hd_decap_3 PHY_84 ();
 scs8hd_decap_3 PHY_85 ();
 scs8hd_tapvpwrvgnd_1 PHY_86 ();
 scs8hd_tapvpwrvgnd_1 PHY_87 ();
 scs8hd_tapvpwrvgnd_1 PHY_88 ();
 scs8hd_tapvpwrvgnd_1 PHY_89 ();
 scs8hd_tapvpwrvgnd_1 PHY_90 ();
 scs8hd_tapvpwrvgnd_1 PHY_91 ();
 scs8hd_tapvpwrvgnd_1 PHY_92 ();
 scs8hd_tapvpwrvgnd_1 PHY_93 ();
 scs8hd_tapvpwrvgnd_1 PHY_94 ();
 scs8hd_tapvpwrvgnd_1 PHY_95 ();
 scs8hd_tapvpwrvgnd_1 PHY_96 ();
 scs8hd_tapvpwrvgnd_1 PHY_97 ();
 scs8hd_tapvpwrvgnd_1 PHY_98 ();
 scs8hd_tapvpwrvgnd_1 PHY_99 ();
 scs8hd_tapvpwrvgnd_1 PHY_100 ();
 scs8hd_tapvpwrvgnd_1 PHY_101 ();
 scs8hd_tapvpwrvgnd_1 PHY_102 ();
 scs8hd_tapvpwrvgnd_1 PHY_103 ();
 scs8hd_tapvpwrvgnd_1 PHY_104 ();
 scs8hd_tapvpwrvgnd_1 PHY_105 ();
 scs8hd_tapvpwrvgnd_1 PHY_106 ();
 scs8hd_tapvpwrvgnd_1 PHY_107 ();
 scs8hd_tapvpwrvgnd_1 PHY_108 ();
 scs8hd_tapvpwrvgnd_1 PHY_109 ();
 scs8hd_tapvpwrvgnd_1 PHY_110 ();
 scs8hd_tapvpwrvgnd_1 PHY_111 ();
 scs8hd_tapvpwrvgnd_1 PHY_112 ();
 scs8hd_tapvpwrvgnd_1 PHY_113 ();
 scs8hd_tapvpwrvgnd_1 PHY_114 ();
 scs8hd_tapvpwrvgnd_1 PHY_115 ();
 scs8hd_tapvpwrvgnd_1 PHY_116 ();
 scs8hd_tapvpwrvgnd_1 PHY_117 ();
 scs8hd_tapvpwrvgnd_1 PHY_118 ();
 scs8hd_tapvpwrvgnd_1 PHY_119 ();
 scs8hd_tapvpwrvgnd_1 PHY_120 ();
 scs8hd_tapvpwrvgnd_1 PHY_121 ();
 scs8hd_tapvpwrvgnd_1 PHY_122 ();
 scs8hd_tapvpwrvgnd_1 PHY_123 ();
 scs8hd_tapvpwrvgnd_1 PHY_124 ();
 scs8hd_tapvpwrvgnd_1 PHY_125 ();
 scs8hd_tapvpwrvgnd_1 PHY_126 ();
 scs8hd_tapvpwrvgnd_1 PHY_127 ();
 scs8hd_tapvpwrvgnd_1 PHY_128 ();
 scs8hd_tapvpwrvgnd_1 PHY_129 ();
 scs8hd_tapvpwrvgnd_1 PHY_130 ();
 scs8hd_tapvpwrvgnd_1 PHY_131 ();
 scs8hd_tapvpwrvgnd_1 PHY_132 ();
 scs8hd_tapvpwrvgnd_1 PHY_133 ();
 scs8hd_tapvpwrvgnd_1 PHY_134 ();
 scs8hd_tapvpwrvgnd_1 PHY_135 ();
 scs8hd_tapvpwrvgnd_1 PHY_136 ();
 scs8hd_tapvpwrvgnd_1 PHY_137 ();
 scs8hd_tapvpwrvgnd_1 PHY_138 ();
 scs8hd_tapvpwrvgnd_1 PHY_139 ();
 scs8hd_tapvpwrvgnd_1 PHY_140 ();
 scs8hd_tapvpwrvgnd_1 PHY_141 ();
 scs8hd_tapvpwrvgnd_1 PHY_142 ();
 scs8hd_tapvpwrvgnd_1 PHY_143 ();
 scs8hd_tapvpwrvgnd_1 PHY_144 ();
 scs8hd_tapvpwrvgnd_1 PHY_145 ();
 scs8hd_tapvpwrvgnd_1 PHY_146 ();
 scs8hd_tapvpwrvgnd_1 PHY_147 ();
 scs8hd_tapvpwrvgnd_1 PHY_148 ();
 scs8hd_tapvpwrvgnd_1 PHY_149 ();
 scs8hd_tapvpwrvgnd_1 PHY_150 ();
 scs8hd_tapvpwrvgnd_1 PHY_151 ();
 scs8hd_tapvpwrvgnd_1 PHY_152 ();
 scs8hd_tapvpwrvgnd_1 PHY_153 ();
 scs8hd_tapvpwrvgnd_1 PHY_154 ();
 scs8hd_tapvpwrvgnd_1 PHY_155 ();
 scs8hd_tapvpwrvgnd_1 PHY_156 ();
 scs8hd_tapvpwrvgnd_1 PHY_157 ();
 scs8hd_tapvpwrvgnd_1 PHY_158 ();
 scs8hd_tapvpwrvgnd_1 PHY_159 ();
 scs8hd_tapvpwrvgnd_1 PHY_160 ();
 scs8hd_tapvpwrvgnd_1 PHY_161 ();
 scs8hd_tapvpwrvgnd_1 PHY_162 ();
 scs8hd_tapvpwrvgnd_1 PHY_163 ();
 scs8hd_tapvpwrvgnd_1 PHY_164 ();
 scs8hd_tapvpwrvgnd_1 PHY_165 ();
 scs8hd_tapvpwrvgnd_1 PHY_166 ();
 scs8hd_tapvpwrvgnd_1 PHY_167 ();
 scs8hd_tapvpwrvgnd_1 PHY_168 ();
 scs8hd_tapvpwrvgnd_1 PHY_169 ();
 scs8hd_tapvpwrvgnd_1 PHY_170 ();
 scs8hd_tapvpwrvgnd_1 PHY_171 ();
 scs8hd_tapvpwrvgnd_1 PHY_172 ();
 scs8hd_tapvpwrvgnd_1 PHY_173 ();
 scs8hd_tapvpwrvgnd_1 PHY_174 ();
 scs8hd_tapvpwrvgnd_1 PHY_175 ();
 scs8hd_tapvpwrvgnd_1 PHY_176 ();
 scs8hd_tapvpwrvgnd_1 PHY_177 ();
 scs8hd_tapvpwrvgnd_1 PHY_178 ();
 scs8hd_tapvpwrvgnd_1 PHY_179 ();
 scs8hd_tapvpwrvgnd_1 PHY_180 ();
 scs8hd_tapvpwrvgnd_1 PHY_181 ();
 scs8hd_tapvpwrvgnd_1 PHY_182 ();
 scs8hd_tapvpwrvgnd_1 PHY_183 ();
 scs8hd_tapvpwrvgnd_1 PHY_184 ();
 scs8hd_tapvpwrvgnd_1 PHY_185 ();
 scs8hd_tapvpwrvgnd_1 PHY_186 ();
 scs8hd_tapvpwrvgnd_1 PHY_187 ();
 scs8hd_tapvpwrvgnd_1 PHY_188 ();
 scs8hd_tapvpwrvgnd_1 PHY_189 ();
 scs8hd_tapvpwrvgnd_1 PHY_190 ();
 scs8hd_tapvpwrvgnd_1 PHY_191 ();
 scs8hd_tapvpwrvgnd_1 PHY_192 ();
 scs8hd_tapvpwrvgnd_1 PHY_193 ();
 scs8hd_tapvpwrvgnd_1 PHY_194 ();
 scs8hd_tapvpwrvgnd_1 PHY_195 ();
 scs8hd_tapvpwrvgnd_1 PHY_196 ();
 scs8hd_tapvpwrvgnd_1 PHY_197 ();
 scs8hd_tapvpwrvgnd_1 PHY_198 ();
 scs8hd_tapvpwrvgnd_1 PHY_199 ();
 scs8hd_tapvpwrvgnd_1 PHY_200 ();
 scs8hd_tapvpwrvgnd_1 PHY_201 ();
 scs8hd_tapvpwrvgnd_1 PHY_202 ();
 scs8hd_tapvpwrvgnd_1 PHY_203 ();
 scs8hd_tapvpwrvgnd_1 PHY_204 ();
 scs8hd_tapvpwrvgnd_1 PHY_205 ();
 scs8hd_tapvpwrvgnd_1 PHY_206 ();
 scs8hd_tapvpwrvgnd_1 PHY_207 ();
 scs8hd_tapvpwrvgnd_1 PHY_208 ();
 scs8hd_tapvpwrvgnd_1 PHY_209 ();
 scs8hd_tapvpwrvgnd_1 PHY_210 ();
 scs8hd_tapvpwrvgnd_1 PHY_211 ();
 scs8hd_tapvpwrvgnd_1 PHY_212 ();
 scs8hd_tapvpwrvgnd_1 PHY_213 ();
 scs8hd_tapvpwrvgnd_1 PHY_214 ();
 scs8hd_tapvpwrvgnd_1 PHY_215 ();
 scs8hd_tapvpwrvgnd_1 PHY_216 ();
 scs8hd_tapvpwrvgnd_1 PHY_217 ();
 scs8hd_tapvpwrvgnd_1 PHY_218 ();
 scs8hd_tapvpwrvgnd_1 PHY_219 ();
 scs8hd_tapvpwrvgnd_1 PHY_220 ();
 scs8hd_tapvpwrvgnd_1 PHY_221 ();
 scs8hd_tapvpwrvgnd_1 PHY_222 ();
 scs8hd_tapvpwrvgnd_1 PHY_223 ();
 scs8hd_tapvpwrvgnd_1 PHY_224 ();
 scs8hd_tapvpwrvgnd_1 PHY_225 ();
 scs8hd_tapvpwrvgnd_1 PHY_226 ();
 scs8hd_tapvpwrvgnd_1 PHY_227 ();
 scs8hd_tapvpwrvgnd_1 PHY_228 ();
 scs8hd_tapvpwrvgnd_1 PHY_229 ();
 scs8hd_tapvpwrvgnd_1 PHY_230 ();
 scs8hd_tapvpwrvgnd_1 PHY_231 ();
 scs8hd_tapvpwrvgnd_1 PHY_232 ();
 scs8hd_tapvpwrvgnd_1 PHY_233 ();
 scs8hd_tapvpwrvgnd_1 PHY_234 ();
 scs8hd_tapvpwrvgnd_1 PHY_235 ();
 scs8hd_tapvpwrvgnd_1 PHY_236 ();
 scs8hd_tapvpwrvgnd_1 PHY_237 ();
 scs8hd_tapvpwrvgnd_1 PHY_238 ();
 scs8hd_tapvpwrvgnd_1 PHY_239 ();
 scs8hd_tapvpwrvgnd_1 PHY_240 ();
 scs8hd_tapvpwrvgnd_1 PHY_241 ();
 scs8hd_tapvpwrvgnd_1 PHY_242 ();
 scs8hd_tapvpwrvgnd_1 PHY_243 ();
 scs8hd_tapvpwrvgnd_1 PHY_244 ();
 scs8hd_tapvpwrvgnd_1 PHY_245 ();
 scs8hd_tapvpwrvgnd_1 PHY_246 ();
 scs8hd_tapvpwrvgnd_1 PHY_247 ();
 scs8hd_tapvpwrvgnd_1 PHY_248 ();
 scs8hd_tapvpwrvgnd_1 PHY_249 ();
 scs8hd_tapvpwrvgnd_1 PHY_250 ();
 scs8hd_tapvpwrvgnd_1 PHY_251 ();
 scs8hd_tapvpwrvgnd_1 PHY_252 ();
 scs8hd_tapvpwrvgnd_1 PHY_253 ();
 scs8hd_tapvpwrvgnd_1 PHY_254 ();
 scs8hd_tapvpwrvgnd_1 PHY_255 ();
 scs8hd_tapvpwrvgnd_1 PHY_256 ();
 scs8hd_tapvpwrvgnd_1 PHY_257 ();
 scs8hd_tapvpwrvgnd_1 PHY_258 ();
 scs8hd_tapvpwrvgnd_1 PHY_259 ();
 scs8hd_tapvpwrvgnd_1 PHY_260 ();
 scs8hd_tapvpwrvgnd_1 PHY_261 ();
 scs8hd_tapvpwrvgnd_1 PHY_262 ();
 scs8hd_tapvpwrvgnd_1 PHY_263 ();
 scs8hd_tapvpwrvgnd_1 PHY_264 ();
 scs8hd_tapvpwrvgnd_1 PHY_265 ();
 scs8hd_diode_2 ANTENNA__CTS_root_A (.DIODE(clk));
 scs8hd_diode_2 ANTENNA__351__A (.DIODE(rst));
 scs8hd_diode_2 ANTENNA__430__B (.DIODE(x[0]));
 scs8hd_diode_2 ANTENNA__504__B (.DIODE(x[10]));
 scs8hd_diode_2 ANTENNA__511__B (.DIODE(x[11]));
 scs8hd_diode_2 ANTENNA__519__B (.DIODE(x[12]));
 scs8hd_diode_2 ANTENNA__526__B (.DIODE(x[13]));
 scs8hd_diode_2 ANTENNA__533__B (.DIODE(x[14]));
 scs8hd_diode_2 ANTENNA__540__B (.DIODE(x[15]));
 scs8hd_diode_2 ANTENNA__547__B (.DIODE(x[16]));
 scs8hd_diode_2 ANTENNA__554__B (.DIODE(x[17]));
 scs8hd_diode_2 ANTENNA__562__B (.DIODE(x[18]));
 scs8hd_diode_2 ANTENNA__569__B (.DIODE(x[19]));
 scs8hd_diode_2 ANTENNA__440__B (.DIODE(x[1]));
 scs8hd_diode_2 ANTENNA__576__B (.DIODE(x[20]));
 scs8hd_diode_2 ANTENNA__583__B (.DIODE(x[21]));
 scs8hd_diode_2 ANTENNA__590__B (.DIODE(x[22]));
 scs8hd_diode_2 ANTENNA__597__B (.DIODE(x[23]));
 scs8hd_diode_2 ANTENNA__605__B (.DIODE(x[24]));
 scs8hd_diode_2 ANTENNA__612__B (.DIODE(x[25]));
 scs8hd_diode_2 ANTENNA__619__B (.DIODE(x[26]));
 scs8hd_diode_2 ANTENNA__626__B (.DIODE(x[27]));
 scs8hd_diode_2 ANTENNA__331__B (.DIODE(x[28]));
 scs8hd_diode_2 ANTENNA__338__B (.DIODE(x[29]));
 scs8hd_diode_2 ANTENNA__447__B (.DIODE(x[2]));
 scs8hd_diode_2 ANTENNA__345__B (.DIODE(x[30]));
 scs8hd_diode_2 ANTENNA__435__B (.DIODE(x[31]));
 scs8hd_diode_2 ANTENNA__454__B (.DIODE(x[3]));
 scs8hd_diode_2 ANTENNA__461__B (.DIODE(x[4]));
 scs8hd_diode_2 ANTENNA__468__B (.DIODE(x[5]));
 scs8hd_diode_2 ANTENNA__476__B (.DIODE(x[6]));
 scs8hd_diode_2 ANTENNA__483__B (.DIODE(x[7]));
 scs8hd_diode_2 ANTENNA__490__B (.DIODE(x[8]));
 scs8hd_diode_2 ANTENNA__497__B (.DIODE(x[9]));
 scs8hd_diode_2 ANTENNA__604__A (.DIODE(y));
 scs8hd_diode_2 ANTENNA__428__A (.DIODE(y));
 scs8hd_diode_2 ANTENNA__655__D (.DIODE(_000_));
 scs8hd_diode_2 ANTENNA__656__D (.DIODE(_001_));
 scs8hd_diode_2 ANTENNA__657__D (.DIODE(_002_));
 scs8hd_diode_2 ANTENNA__658__D (.DIODE(_003_));
 scs8hd_diode_2 ANTENNA__659__D (.DIODE(_004_));
 scs8hd_diode_2 ANTENNA__660__D (.DIODE(_005_));
 scs8hd_diode_2 ANTENNA__661__D (.DIODE(_006_));
 scs8hd_diode_2 ANTENNA__662__D (.DIODE(_007_));
 scs8hd_diode_2 ANTENNA__663__D (.DIODE(_008_));
 scs8hd_diode_2 ANTENNA__664__D (.DIODE(_009_));
 scs8hd_diode_2 ANTENNA__665__D (.DIODE(_010_));
 scs8hd_diode_2 ANTENNA__666__D (.DIODE(_011_));
 scs8hd_diode_2 ANTENNA__667__D (.DIODE(_012_));
 scs8hd_diode_2 ANTENNA__668__D (.DIODE(_013_));
 scs8hd_diode_2 ANTENNA__669__D (.DIODE(_014_));
 scs8hd_diode_2 ANTENNA__670__D (.DIODE(_015_));
 scs8hd_diode_2 ANTENNA__671__D (.DIODE(_016_));
 scs8hd_diode_2 ANTENNA__672__D (.DIODE(_017_));
 scs8hd_diode_2 ANTENNA__673__D (.DIODE(_018_));
 scs8hd_diode_2 ANTENNA__674__D (.DIODE(_019_));
 scs8hd_diode_2 ANTENNA__637__D (.DIODE(_020_));
 scs8hd_diode_2 ANTENNA__638__D (.DIODE(_021_));
 scs8hd_diode_2 ANTENNA__675__D (.DIODE(_022_));
 scs8hd_diode_2 ANTENNA__676__D (.DIODE(_023_));
 scs8hd_diode_2 ANTENNA__677__D (.DIODE(_024_));
 scs8hd_diode_2 ANTENNA__678__D (.DIODE(_025_));
 scs8hd_diode_2 ANTENNA__679__D (.DIODE(_026_));
 scs8hd_diode_2 ANTENNA__680__D (.DIODE(_027_));
 scs8hd_diode_2 ANTENNA__681__D (.DIODE(_028_));
 scs8hd_diode_2 ANTENNA__682__D (.DIODE(_029_));
 scs8hd_diode_2 ANTENNA__683__D (.DIODE(_030_));
 scs8hd_diode_2 ANTENNA__684__D (.DIODE(_031_));
 scs8hd_diode_2 ANTENNA__685__D (.DIODE(_032_));
 scs8hd_diode_2 ANTENNA__686__D (.DIODE(_033_));
 scs8hd_diode_2 ANTENNA__687__D (.DIODE(_034_));
 scs8hd_diode_2 ANTENNA__688__D (.DIODE(_035_));
 scs8hd_diode_2 ANTENNA__689__D (.DIODE(_036_));
 scs8hd_diode_2 ANTENNA__690__D (.DIODE(_037_));
 scs8hd_diode_2 ANTENNA__691__D (.DIODE(_038_));
 scs8hd_diode_2 ANTENNA__692__D (.DIODE(_039_));
 scs8hd_diode_2 ANTENNA__693__D (.DIODE(_040_));
 scs8hd_diode_2 ANTENNA__694__D (.DIODE(_041_));
 scs8hd_diode_2 ANTENNA__639__D (.DIODE(_042_));
 scs8hd_diode_2 ANTENNA__640__D (.DIODE(_043_));
 scs8hd_diode_2 ANTENNA__695__D (.DIODE(_044_));
 scs8hd_diode_2 ANTENNA__696__D (.DIODE(_045_));
 scs8hd_diode_2 ANTENNA__641__D (.DIODE(_046_));
 scs8hd_diode_2 ANTENNA__642__D (.DIODE(_047_));
 scs8hd_diode_2 ANTENNA__643__D (.DIODE(_048_));
 scs8hd_diode_2 ANTENNA__644__D (.DIODE(_049_));
 scs8hd_diode_2 ANTENNA__645__D (.DIODE(_050_));
 scs8hd_diode_2 ANTENNA__646__D (.DIODE(_051_));
 scs8hd_diode_2 ANTENNA__647__D (.DIODE(_052_));
 scs8hd_diode_2 ANTENNA__648__D (.DIODE(_053_));
 scs8hd_diode_2 ANTENNA__649__D (.DIODE(_054_));
 scs8hd_diode_2 ANTENNA__650__D (.DIODE(_055_));
 scs8hd_diode_2 ANTENNA__651__D (.DIODE(_056_));
 scs8hd_diode_2 ANTENNA__652__D (.DIODE(_057_));
 scs8hd_diode_2 ANTENNA__653__D (.DIODE(_058_));
 scs8hd_diode_2 ANTENNA__654__D (.DIODE(_059_));
 scs8hd_diode_2 ANTENNA__633__D (.DIODE(_060_));
 scs8hd_diode_2 ANTENNA__636__D (.DIODE(_061_));
 scs8hd_diode_2 ANTENNA__635__D (.DIODE(_062_));
 scs8hd_diode_2 ANTENNA__437__B1N (.DIODE(_062_));
 scs8hd_diode_2 ANTENNA__506__B1 (.DIODE(_063_));
 scs8hd_diode_2 ANTENNA__502__A (.DIODE(_063_));
 scs8hd_diode_2 ANTENNA__513__B1 (.DIODE(_064_));
 scs8hd_diode_2 ANTENNA__509__A (.DIODE(_064_));
 scs8hd_diode_2 ANTENNA__521__B1 (.DIODE(_065_));
 scs8hd_diode_2 ANTENNA__516__A (.DIODE(_065_));
 scs8hd_diode_2 ANTENNA__528__B1 (.DIODE(_066_));
 scs8hd_diode_2 ANTENNA__524__A (.DIODE(_066_));
 scs8hd_diode_2 ANTENNA__535__B1 (.DIODE(_067_));
 scs8hd_diode_2 ANTENNA__531__A (.DIODE(_067_));
 scs8hd_diode_2 ANTENNA__542__B1 (.DIODE(_068_));
 scs8hd_diode_2 ANTENNA__538__A (.DIODE(_068_));
 scs8hd_diode_2 ANTENNA__549__B1 (.DIODE(_069_));
 scs8hd_diode_2 ANTENNA__545__A (.DIODE(_069_));
 scs8hd_diode_2 ANTENNA__556__B1 (.DIODE(_070_));
 scs8hd_diode_2 ANTENNA__552__A (.DIODE(_070_));
 scs8hd_diode_2 ANTENNA__564__B1 (.DIODE(_071_));
 scs8hd_diode_2 ANTENNA__559__A (.DIODE(_071_));
 scs8hd_diode_2 ANTENNA__571__B1 (.DIODE(_072_));
 scs8hd_diode_2 ANTENNA__567__A (.DIODE(_072_));
 scs8hd_diode_2 ANTENNA__442__B1 (.DIODE(_073_));
 scs8hd_diode_2 ANTENNA__438__A (.DIODE(_073_));
 scs8hd_diode_2 ANTENNA__578__B1 (.DIODE(_074_));
 scs8hd_diode_2 ANTENNA__574__A (.DIODE(_074_));
 scs8hd_diode_2 ANTENNA__585__B1 (.DIODE(_075_));
 scs8hd_diode_2 ANTENNA__581__A (.DIODE(_075_));
 scs8hd_diode_2 ANTENNA__592__B1 (.DIODE(_076_));
 scs8hd_diode_2 ANTENNA__588__A (.DIODE(_076_));
 scs8hd_diode_2 ANTENNA__599__B1 (.DIODE(_077_));
 scs8hd_diode_2 ANTENNA__595__A (.DIODE(_077_));
 scs8hd_diode_2 ANTENNA__607__B1 (.DIODE(_078_));
 scs8hd_diode_2 ANTENNA__602__A (.DIODE(_078_));
 scs8hd_diode_2 ANTENNA__614__B1 (.DIODE(_079_));
 scs8hd_diode_2 ANTENNA__610__A (.DIODE(_079_));
 scs8hd_diode_2 ANTENNA__621__B1 (.DIODE(_080_));
 scs8hd_diode_2 ANTENNA__617__A (.DIODE(_080_));
 scs8hd_diode_2 ANTENNA__628__B1 (.DIODE(_081_));
 scs8hd_diode_2 ANTENNA__624__A (.DIODE(_081_));
 scs8hd_diode_2 ANTENNA__631__A (.DIODE(_082_));
 scs8hd_diode_2 ANTENNA__333__B1 (.DIODE(_082_));
 scs8hd_diode_2 ANTENNA__340__B1 (.DIODE(_083_));
 scs8hd_diode_2 ANTENNA__336__A (.DIODE(_083_));
 scs8hd_diode_2 ANTENNA__449__B1 (.DIODE(_084_));
 scs8hd_diode_2 ANTENNA__445__A (.DIODE(_084_));
 scs8hd_diode_2 ANTENNA__347__B1 (.DIODE(_085_));
 scs8hd_diode_2 ANTENNA__343__A (.DIODE(_085_));
 scs8hd_diode_2 ANTENNA__456__B1 (.DIODE(_086_));
 scs8hd_diode_2 ANTENNA__452__A (.DIODE(_086_));
 scs8hd_diode_2 ANTENNA__463__B1 (.DIODE(_087_));
 scs8hd_diode_2 ANTENNA__459__A (.DIODE(_087_));
 scs8hd_diode_2 ANTENNA__470__B1 (.DIODE(_088_));
 scs8hd_diode_2 ANTENNA__466__A (.DIODE(_088_));
 scs8hd_diode_2 ANTENNA__478__B1 (.DIODE(_089_));
 scs8hd_diode_2 ANTENNA__473__A (.DIODE(_089_));
 scs8hd_diode_2 ANTENNA__485__B1 (.DIODE(_090_));
 scs8hd_diode_2 ANTENNA__481__A (.DIODE(_090_));
 scs8hd_diode_2 ANTENNA__492__B1 (.DIODE(_091_));
 scs8hd_diode_2 ANTENNA__488__A (.DIODE(_091_));
 scs8hd_diode_2 ANTENNA__499__B1 (.DIODE(_092_));
 scs8hd_diode_2 ANTENNA__495__A (.DIODE(_092_));
 scs8hd_diode_2 ANTENNA__633__RESETB (.DIODE(_093_));
 scs8hd_diode_2 ANTENNA__634__RESETB (.DIODE(_094_));
 scs8hd_diode_2 ANTENNA__635__RESETB (.DIODE(_095_));
 scs8hd_diode_2 ANTENNA__636__RESETB (.DIODE(_096_));
 scs8hd_diode_2 ANTENNA__637__RESETB (.DIODE(_097_));
 scs8hd_diode_2 ANTENNA__638__RESETB (.DIODE(_098_));
 scs8hd_diode_2 ANTENNA__639__RESETB (.DIODE(_099_));
 scs8hd_diode_2 ANTENNA__640__RESETB (.DIODE(_100_));
 scs8hd_diode_2 ANTENNA__641__RESETB (.DIODE(_101_));
 scs8hd_diode_2 ANTENNA__642__RESETB (.DIODE(_102_));
 scs8hd_diode_2 ANTENNA__643__RESETB (.DIODE(_103_));
 scs8hd_diode_2 ANTENNA__644__RESETB (.DIODE(_104_));
 scs8hd_diode_2 ANTENNA__645__RESETB (.DIODE(_105_));
 scs8hd_diode_2 ANTENNA__646__RESETB (.DIODE(_106_));
 scs8hd_diode_2 ANTENNA__647__RESETB (.DIODE(_107_));
 scs8hd_diode_2 ANTENNA__648__RESETB (.DIODE(_108_));
 scs8hd_diode_2 ANTENNA__649__RESETB (.DIODE(_109_));
 scs8hd_diode_2 ANTENNA__650__RESETB (.DIODE(_110_));
 scs8hd_diode_2 ANTENNA__651__RESETB (.DIODE(_111_));
 scs8hd_diode_2 ANTENNA__652__RESETB (.DIODE(_112_));
 scs8hd_diode_2 ANTENNA__653__RESETB (.DIODE(_113_));
 scs8hd_diode_2 ANTENNA__654__RESETB (.DIODE(_114_));
 scs8hd_diode_2 ANTENNA__655__RESETB (.DIODE(_115_));
 scs8hd_diode_2 ANTENNA__656__RESETB (.DIODE(_116_));
 scs8hd_diode_2 ANTENNA__657__RESETB (.DIODE(_117_));
 scs8hd_diode_2 ANTENNA__658__RESETB (.DIODE(_118_));
 scs8hd_diode_2 ANTENNA__659__RESETB (.DIODE(_119_));
 scs8hd_diode_2 ANTENNA__660__RESETB (.DIODE(_120_));
 scs8hd_diode_2 ANTENNA__661__RESETB (.DIODE(_121_));
 scs8hd_diode_2 ANTENNA__662__RESETB (.DIODE(_122_));
 scs8hd_diode_2 ANTENNA__663__RESETB (.DIODE(_123_));
 scs8hd_diode_2 ANTENNA__664__RESETB (.DIODE(_124_));
 scs8hd_diode_2 ANTENNA__665__RESETB (.DIODE(_125_));
 scs8hd_diode_2 ANTENNA__666__RESETB (.DIODE(_126_));
 scs8hd_diode_2 ANTENNA__667__RESETB (.DIODE(_127_));
 scs8hd_diode_2 ANTENNA__668__RESETB (.DIODE(_128_));
 scs8hd_diode_2 ANTENNA__669__RESETB (.DIODE(_129_));
 scs8hd_diode_2 ANTENNA__670__RESETB (.DIODE(_130_));
 scs8hd_diode_2 ANTENNA__671__RESETB (.DIODE(_131_));
 scs8hd_diode_2 ANTENNA__672__RESETB (.DIODE(_132_));
 scs8hd_diode_2 ANTENNA__673__RESETB (.DIODE(_133_));
 scs8hd_diode_2 ANTENNA__674__RESETB (.DIODE(_134_));
 scs8hd_diode_2 ANTENNA__675__RESETB (.DIODE(_135_));
 scs8hd_diode_2 ANTENNA__676__RESETB (.DIODE(_136_));
 scs8hd_diode_2 ANTENNA__677__RESETB (.DIODE(_137_));
 scs8hd_diode_2 ANTENNA__678__RESETB (.DIODE(_138_));
 scs8hd_diode_2 ANTENNA__679__RESETB (.DIODE(_139_));
 scs8hd_diode_2 ANTENNA__680__RESETB (.DIODE(_140_));
 scs8hd_diode_2 ANTENNA__681__RESETB (.DIODE(_141_));
 scs8hd_diode_2 ANTENNA__682__RESETB (.DIODE(_142_));
 scs8hd_diode_2 ANTENNA__683__RESETB (.DIODE(_143_));
 scs8hd_diode_2 ANTENNA__684__RESETB (.DIODE(_144_));
 scs8hd_diode_2 ANTENNA__685__RESETB (.DIODE(_145_));
 scs8hd_diode_2 ANTENNA__686__RESETB (.DIODE(_146_));
 scs8hd_diode_2 ANTENNA__687__RESETB (.DIODE(_147_));
 scs8hd_diode_2 ANTENNA__688__RESETB (.DIODE(_148_));
 scs8hd_diode_2 ANTENNA__689__RESETB (.DIODE(_149_));
 scs8hd_diode_2 ANTENNA__690__RESETB (.DIODE(_150_));
 scs8hd_diode_2 ANTENNA__691__RESETB (.DIODE(_151_));
 scs8hd_diode_2 ANTENNA__692__RESETB (.DIODE(_152_));
 scs8hd_diode_2 ANTENNA__693__RESETB (.DIODE(_153_));
 scs8hd_diode_2 ANTENNA__694__RESETB (.DIODE(_154_));
 scs8hd_diode_2 ANTENNA__695__RESETB (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__357__A (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__356__A (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__355__A (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__354__A (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__353__A (.DIODE(_155_));
 scs8hd_diode_2 ANTENNA__696__RESETB (.DIODE(_156_));
 scs8hd_diode_2 ANTENNA__416__A (.DIODE(_157_));
 scs8hd_diode_2 ANTENNA__373__A (.DIODE(_157_));
 scs8hd_diode_2 ANTENNA__358__A (.DIODE(_157_));
 scs8hd_diode_2 ANTENNA__352__A (.DIODE(_157_));
 scs8hd_diode_2 ANTENNA__425__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__424__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__423__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__366__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__359__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__350__A (.DIODE(_158_));
 scs8hd_diode_2 ANTENNA__365__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__364__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__363__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__362__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__361__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__360__A (.DIODE(_159_));
 scs8hd_diode_2 ANTENNA__372__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__371__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__370__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__369__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__368__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__367__A (.DIODE(_160_));
 scs8hd_diode_2 ANTENNA__409__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__402__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__395__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__388__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__381__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__374__A (.DIODE(_161_));
 scs8hd_diode_2 ANTENNA__380__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__379__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__378__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__377__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__376__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__375__A (.DIODE(_162_));
 scs8hd_diode_2 ANTENNA__387__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__386__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__385__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__384__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__383__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__382__A (.DIODE(_163_));
 scs8hd_diode_2 ANTENNA__394__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__393__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__392__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__391__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__390__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__389__A (.DIODE(_164_));
 scs8hd_diode_2 ANTENNA__401__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__400__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__399__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__398__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__397__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__396__A (.DIODE(_165_));
 scs8hd_diode_2 ANTENNA__408__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__407__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__406__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__405__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__404__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__403__A (.DIODE(_166_));
 scs8hd_diode_2 ANTENNA__415__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__414__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__413__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__412__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__411__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__410__A (.DIODE(_167_));
 scs8hd_diode_2 ANTENNA__422__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__421__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__420__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__419__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__418__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__417__A (.DIODE(_168_));
 scs8hd_diode_2 ANTENNA__433__A1N (.DIODE(_169_));
 scs8hd_diode_2 ANTENNA__432__A1 (.DIODE(_169_));
 scs8hd_diode_2 ANTENNA__433__A2N (.DIODE(_170_));
 scs8hd_diode_2 ANTENNA__432__A2 (.DIODE(_170_));
 scs8hd_diode_2 ANTENNA__561__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__518__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__475__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__435__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__429__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__345__A (.DIODE(_171_));
 scs8hd_diode_2 ANTENNA__468__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__461__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__454__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__447__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__440__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__430__A (.DIODE(_172_));
 scs8hd_diode_2 ANTENNA__431__A (.DIODE(_173_));
 scs8hd_diode_2 ANTENNA__434__A (.DIODE(_174_));
 scs8hd_diode_2 ANTENNA__433__B1 (.DIODE(_174_));
 scs8hd_diode_2 ANTENNA__434__B (.DIODE(_175_));
 scs8hd_diode_2 ANTENNA__433__B2 (.DIODE(_175_));
 scs8hd_diode_2 ANTENNA__437__A2 (.DIODE(_176_));
 scs8hd_diode_2 ANTENNA__436__B (.DIODE(_176_));
 scs8hd_diode_2 ANTENNA__443__A1N (.DIODE(_177_));
 scs8hd_diode_2 ANTENNA__442__A1 (.DIODE(_177_));
 scs8hd_diode_2 ANTENNA__443__A2N (.DIODE(_178_));
 scs8hd_diode_2 ANTENNA__442__A2 (.DIODE(_178_));
 scs8hd_diode_2 ANTENNA__441__A (.DIODE(_179_));
 scs8hd_diode_2 ANTENNA__444__A (.DIODE(_180_));
 scs8hd_diode_2 ANTENNA__443__B1 (.DIODE(_180_));
 scs8hd_diode_2 ANTENNA__444__B (.DIODE(_181_));
 scs8hd_diode_2 ANTENNA__443__B2 (.DIODE(_181_));
 scs8hd_diode_2 ANTENNA__450__A1N (.DIODE(_182_));
 scs8hd_diode_2 ANTENNA__449__A1 (.DIODE(_182_));
 scs8hd_diode_2 ANTENNA__450__A2N (.DIODE(_183_));
 scs8hd_diode_2 ANTENNA__449__A2 (.DIODE(_183_));
 scs8hd_diode_2 ANTENNA__448__A (.DIODE(_184_));
 scs8hd_diode_2 ANTENNA__451__A (.DIODE(_185_));
 scs8hd_diode_2 ANTENNA__450__B1 (.DIODE(_185_));
 scs8hd_diode_2 ANTENNA__451__B (.DIODE(_186_));
 scs8hd_diode_2 ANTENNA__450__B2 (.DIODE(_186_));
 scs8hd_diode_2 ANTENNA__457__A1N (.DIODE(_187_));
 scs8hd_diode_2 ANTENNA__456__A1 (.DIODE(_187_));
 scs8hd_diode_2 ANTENNA__457__A2N (.DIODE(_188_));
 scs8hd_diode_2 ANTENNA__456__A2 (.DIODE(_188_));
 scs8hd_diode_2 ANTENNA__455__A (.DIODE(_189_));
 scs8hd_diode_2 ANTENNA__458__A (.DIODE(_190_));
 scs8hd_diode_2 ANTENNA__457__B1 (.DIODE(_190_));
 scs8hd_diode_2 ANTENNA__458__B (.DIODE(_191_));
 scs8hd_diode_2 ANTENNA__457__B2 (.DIODE(_191_));
 scs8hd_diode_2 ANTENNA__464__A1N (.DIODE(_192_));
 scs8hd_diode_2 ANTENNA__463__A1 (.DIODE(_192_));
 scs8hd_diode_2 ANTENNA__464__A2N (.DIODE(_193_));
 scs8hd_diode_2 ANTENNA__463__A2 (.DIODE(_193_));
 scs8hd_diode_2 ANTENNA__462__A (.DIODE(_194_));
 scs8hd_diode_2 ANTENNA__465__A (.DIODE(_195_));
 scs8hd_diode_2 ANTENNA__464__B1 (.DIODE(_195_));
 scs8hd_diode_2 ANTENNA__465__B (.DIODE(_196_));
 scs8hd_diode_2 ANTENNA__464__B2 (.DIODE(_196_));
 scs8hd_diode_2 ANTENNA__471__A1N (.DIODE(_197_));
 scs8hd_diode_2 ANTENNA__470__A1 (.DIODE(_197_));
 scs8hd_diode_2 ANTENNA__471__A2N (.DIODE(_198_));
 scs8hd_diode_2 ANTENNA__470__A2 (.DIODE(_198_));
 scs8hd_diode_2 ANTENNA__469__A (.DIODE(_199_));
 scs8hd_diode_2 ANTENNA__472__A (.DIODE(_200_));
 scs8hd_diode_2 ANTENNA__471__B1 (.DIODE(_200_));
 scs8hd_diode_2 ANTENNA__472__B (.DIODE(_201_));
 scs8hd_diode_2 ANTENNA__471__B2 (.DIODE(_201_));
 scs8hd_diode_2 ANTENNA__479__A1N (.DIODE(_202_));
 scs8hd_diode_2 ANTENNA__478__A1 (.DIODE(_202_));
 scs8hd_diode_2 ANTENNA__479__A2N (.DIODE(_203_));
 scs8hd_diode_2 ANTENNA__478__A2 (.DIODE(_203_));
 scs8hd_diode_2 ANTENNA__511__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__504__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__497__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__490__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__483__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__476__A (.DIODE(_204_));
 scs8hd_diode_2 ANTENNA__477__A (.DIODE(_205_));
 scs8hd_diode_2 ANTENNA__480__A (.DIODE(_206_));
 scs8hd_diode_2 ANTENNA__479__B1 (.DIODE(_206_));
 scs8hd_diode_2 ANTENNA__480__B (.DIODE(_207_));
 scs8hd_diode_2 ANTENNA__479__B2 (.DIODE(_207_));
 scs8hd_diode_2 ANTENNA__486__A1N (.DIODE(_208_));
 scs8hd_diode_2 ANTENNA__485__A1 (.DIODE(_208_));
 scs8hd_diode_2 ANTENNA__486__A2N (.DIODE(_209_));
 scs8hd_diode_2 ANTENNA__485__A2 (.DIODE(_209_));
 scs8hd_diode_2 ANTENNA__484__A (.DIODE(_210_));
 scs8hd_diode_2 ANTENNA__487__A (.DIODE(_211_));
 scs8hd_diode_2 ANTENNA__486__B1 (.DIODE(_211_));
 scs8hd_diode_2 ANTENNA__487__B (.DIODE(_212_));
 scs8hd_diode_2 ANTENNA__486__B2 (.DIODE(_212_));
 scs8hd_diode_2 ANTENNA__493__A1N (.DIODE(_213_));
 scs8hd_diode_2 ANTENNA__492__A1 (.DIODE(_213_));
 scs8hd_diode_2 ANTENNA__493__A2N (.DIODE(_214_));
 scs8hd_diode_2 ANTENNA__492__A2 (.DIODE(_214_));
 scs8hd_diode_2 ANTENNA__491__A (.DIODE(_215_));
 scs8hd_diode_2 ANTENNA__494__A (.DIODE(_216_));
 scs8hd_diode_2 ANTENNA__493__B1 (.DIODE(_216_));
 scs8hd_diode_2 ANTENNA__494__B (.DIODE(_217_));
 scs8hd_diode_2 ANTENNA__493__B2 (.DIODE(_217_));
 scs8hd_diode_2 ANTENNA__500__A1N (.DIODE(_218_));
 scs8hd_diode_2 ANTENNA__499__A1 (.DIODE(_218_));
 scs8hd_diode_2 ANTENNA__500__A2N (.DIODE(_219_));
 scs8hd_diode_2 ANTENNA__499__A2 (.DIODE(_219_));
 scs8hd_diode_2 ANTENNA__498__A (.DIODE(_220_));
 scs8hd_diode_2 ANTENNA__501__A (.DIODE(_221_));
 scs8hd_diode_2 ANTENNA__500__B1 (.DIODE(_221_));
 scs8hd_diode_2 ANTENNA__501__B (.DIODE(_222_));
 scs8hd_diode_2 ANTENNA__500__B2 (.DIODE(_222_));
 scs8hd_diode_2 ANTENNA__507__A1N (.DIODE(_223_));
 scs8hd_diode_2 ANTENNA__506__A1 (.DIODE(_223_));
 scs8hd_diode_2 ANTENNA__507__A2N (.DIODE(_224_));
 scs8hd_diode_2 ANTENNA__506__A2 (.DIODE(_224_));
 scs8hd_diode_2 ANTENNA__505__A (.DIODE(_225_));
 scs8hd_diode_2 ANTENNA__508__A (.DIODE(_226_));
 scs8hd_diode_2 ANTENNA__507__B1 (.DIODE(_226_));
 scs8hd_diode_2 ANTENNA__508__B (.DIODE(_227_));
 scs8hd_diode_2 ANTENNA__507__B2 (.DIODE(_227_));
 scs8hd_diode_2 ANTENNA__514__A1N (.DIODE(_228_));
 scs8hd_diode_2 ANTENNA__513__A1 (.DIODE(_228_));
 scs8hd_diode_2 ANTENNA__514__A2N (.DIODE(_229_));
 scs8hd_diode_2 ANTENNA__513__A2 (.DIODE(_229_));
 scs8hd_diode_2 ANTENNA__512__A (.DIODE(_230_));
 scs8hd_diode_2 ANTENNA__515__A (.DIODE(_231_));
 scs8hd_diode_2 ANTENNA__514__B1 (.DIODE(_231_));
 scs8hd_diode_2 ANTENNA__515__B (.DIODE(_232_));
 scs8hd_diode_2 ANTENNA__514__B2 (.DIODE(_232_));
 scs8hd_diode_2 ANTENNA__522__A1N (.DIODE(_233_));
 scs8hd_diode_2 ANTENNA__521__A1 (.DIODE(_233_));
 scs8hd_diode_2 ANTENNA__522__A2N (.DIODE(_234_));
 scs8hd_diode_2 ANTENNA__521__A2 (.DIODE(_234_));
 scs8hd_diode_2 ANTENNA__554__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__547__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__540__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__533__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__526__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__519__A (.DIODE(_235_));
 scs8hd_diode_2 ANTENNA__520__A (.DIODE(_236_));
 scs8hd_diode_2 ANTENNA__523__A (.DIODE(_237_));
 scs8hd_diode_2 ANTENNA__522__B1 (.DIODE(_237_));
 scs8hd_diode_2 ANTENNA__523__B (.DIODE(_238_));
 scs8hd_diode_2 ANTENNA__522__B2 (.DIODE(_238_));
 scs8hd_diode_2 ANTENNA__529__A1N (.DIODE(_239_));
 scs8hd_diode_2 ANTENNA__528__A1 (.DIODE(_239_));
 scs8hd_diode_2 ANTENNA__529__A2N (.DIODE(_240_));
 scs8hd_diode_2 ANTENNA__528__A2 (.DIODE(_240_));
 scs8hd_diode_2 ANTENNA__527__A (.DIODE(_241_));
 scs8hd_diode_2 ANTENNA__530__A (.DIODE(_242_));
 scs8hd_diode_2 ANTENNA__529__B1 (.DIODE(_242_));
 scs8hd_diode_2 ANTENNA__530__B (.DIODE(_243_));
 scs8hd_diode_2 ANTENNA__529__B2 (.DIODE(_243_));
 scs8hd_diode_2 ANTENNA__536__A1N (.DIODE(_244_));
 scs8hd_diode_2 ANTENNA__535__A1 (.DIODE(_244_));
 scs8hd_diode_2 ANTENNA__536__A2N (.DIODE(_245_));
 scs8hd_diode_2 ANTENNA__535__A2 (.DIODE(_245_));
 scs8hd_diode_2 ANTENNA__534__A (.DIODE(_246_));
 scs8hd_diode_2 ANTENNA__537__A (.DIODE(_247_));
 scs8hd_diode_2 ANTENNA__536__B1 (.DIODE(_247_));
 scs8hd_diode_2 ANTENNA__537__B (.DIODE(_248_));
 scs8hd_diode_2 ANTENNA__536__B2 (.DIODE(_248_));
 scs8hd_diode_2 ANTENNA__543__A1N (.DIODE(_249_));
 scs8hd_diode_2 ANTENNA__542__A1 (.DIODE(_249_));
 scs8hd_diode_2 ANTENNA__543__A2N (.DIODE(_250_));
 scs8hd_diode_2 ANTENNA__542__A2 (.DIODE(_250_));
 scs8hd_diode_2 ANTENNA__541__A (.DIODE(_251_));
 scs8hd_diode_2 ANTENNA__544__A (.DIODE(_252_));
 scs8hd_diode_2 ANTENNA__543__B1 (.DIODE(_252_));
 scs8hd_diode_2 ANTENNA__544__B (.DIODE(_253_));
 scs8hd_diode_2 ANTENNA__543__B2 (.DIODE(_253_));
 scs8hd_diode_2 ANTENNA__550__A1N (.DIODE(_254_));
 scs8hd_diode_2 ANTENNA__549__A1 (.DIODE(_254_));
 scs8hd_diode_2 ANTENNA__550__A2N (.DIODE(_255_));
 scs8hd_diode_2 ANTENNA__549__A2 (.DIODE(_255_));
 scs8hd_diode_2 ANTENNA__548__A (.DIODE(_256_));
 scs8hd_diode_2 ANTENNA__551__A (.DIODE(_257_));
 scs8hd_diode_2 ANTENNA__550__B1 (.DIODE(_257_));
 scs8hd_diode_2 ANTENNA__551__B (.DIODE(_258_));
 scs8hd_diode_2 ANTENNA__550__B2 (.DIODE(_258_));
 scs8hd_diode_2 ANTENNA__557__A1N (.DIODE(_259_));
 scs8hd_diode_2 ANTENNA__556__A1 (.DIODE(_259_));
 scs8hd_diode_2 ANTENNA__557__A2N (.DIODE(_260_));
 scs8hd_diode_2 ANTENNA__556__A2 (.DIODE(_260_));
 scs8hd_diode_2 ANTENNA__555__A (.DIODE(_261_));
 scs8hd_diode_2 ANTENNA__558__A (.DIODE(_262_));
 scs8hd_diode_2 ANTENNA__557__B1 (.DIODE(_262_));
 scs8hd_diode_2 ANTENNA__558__B (.DIODE(_263_));
 scs8hd_diode_2 ANTENNA__557__B2 (.DIODE(_263_));
 scs8hd_diode_2 ANTENNA__565__A1N (.DIODE(_264_));
 scs8hd_diode_2 ANTENNA__564__A1 (.DIODE(_264_));
 scs8hd_diode_2 ANTENNA__565__A2N (.DIODE(_265_));
 scs8hd_diode_2 ANTENNA__564__A2 (.DIODE(_265_));
 scs8hd_diode_2 ANTENNA__597__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__590__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__583__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__576__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__569__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__562__A (.DIODE(_266_));
 scs8hd_diode_2 ANTENNA__563__A (.DIODE(_267_));
 scs8hd_diode_2 ANTENNA__566__A (.DIODE(_268_));
 scs8hd_diode_2 ANTENNA__565__B1 (.DIODE(_268_));
 scs8hd_diode_2 ANTENNA__566__B (.DIODE(_269_));
 scs8hd_diode_2 ANTENNA__565__B2 (.DIODE(_269_));
 scs8hd_diode_2 ANTENNA__572__A1N (.DIODE(_270_));
 scs8hd_diode_2 ANTENNA__571__A1 (.DIODE(_270_));
 scs8hd_diode_2 ANTENNA__572__A2N (.DIODE(_271_));
 scs8hd_diode_2 ANTENNA__571__A2 (.DIODE(_271_));
 scs8hd_diode_2 ANTENNA__570__A (.DIODE(_272_));
 scs8hd_diode_2 ANTENNA__573__A (.DIODE(_273_));
 scs8hd_diode_2 ANTENNA__572__B1 (.DIODE(_273_));
 scs8hd_diode_2 ANTENNA__573__B (.DIODE(_274_));
 scs8hd_diode_2 ANTENNA__572__B2 (.DIODE(_274_));
 scs8hd_diode_2 ANTENNA__579__A1N (.DIODE(_275_));
 scs8hd_diode_2 ANTENNA__578__A1 (.DIODE(_275_));
 scs8hd_diode_2 ANTENNA__579__A2N (.DIODE(_276_));
 scs8hd_diode_2 ANTENNA__578__A2 (.DIODE(_276_));
 scs8hd_diode_2 ANTENNA__577__A (.DIODE(_277_));
 scs8hd_diode_2 ANTENNA__580__A (.DIODE(_278_));
 scs8hd_diode_2 ANTENNA__579__B1 (.DIODE(_278_));
 scs8hd_diode_2 ANTENNA__580__B (.DIODE(_279_));
 scs8hd_diode_2 ANTENNA__579__B2 (.DIODE(_279_));
 scs8hd_diode_2 ANTENNA__586__A1N (.DIODE(_280_));
 scs8hd_diode_2 ANTENNA__585__A1 (.DIODE(_280_));
 scs8hd_diode_2 ANTENNA__586__A2N (.DIODE(_281_));
 scs8hd_diode_2 ANTENNA__585__A2 (.DIODE(_281_));
 scs8hd_diode_2 ANTENNA__584__A (.DIODE(_282_));
 scs8hd_diode_2 ANTENNA__587__A (.DIODE(_283_));
 scs8hd_diode_2 ANTENNA__586__B1 (.DIODE(_283_));
 scs8hd_diode_2 ANTENNA__587__B (.DIODE(_284_));
 scs8hd_diode_2 ANTENNA__586__B2 (.DIODE(_284_));
 scs8hd_diode_2 ANTENNA__593__A1N (.DIODE(_285_));
 scs8hd_diode_2 ANTENNA__592__A1 (.DIODE(_285_));
 scs8hd_diode_2 ANTENNA__593__A2N (.DIODE(_286_));
 scs8hd_diode_2 ANTENNA__592__A2 (.DIODE(_286_));
 scs8hd_diode_2 ANTENNA__591__A (.DIODE(_287_));
 scs8hd_diode_2 ANTENNA__594__A (.DIODE(_288_));
 scs8hd_diode_2 ANTENNA__593__B1 (.DIODE(_288_));
 scs8hd_diode_2 ANTENNA__594__B (.DIODE(_289_));
 scs8hd_diode_2 ANTENNA__593__B2 (.DIODE(_289_));
 scs8hd_diode_2 ANTENNA__600__A1N (.DIODE(_290_));
 scs8hd_diode_2 ANTENNA__599__A1 (.DIODE(_290_));
 scs8hd_diode_2 ANTENNA__600__A2N (.DIODE(_291_));
 scs8hd_diode_2 ANTENNA__599__A2 (.DIODE(_291_));
 scs8hd_diode_2 ANTENNA__598__A (.DIODE(_292_));
 scs8hd_diode_2 ANTENNA__601__A (.DIODE(_293_));
 scs8hd_diode_2 ANTENNA__600__B1 (.DIODE(_293_));
 scs8hd_diode_2 ANTENNA__601__B (.DIODE(_294_));
 scs8hd_diode_2 ANTENNA__600__B2 (.DIODE(_294_));
 scs8hd_diode_2 ANTENNA__608__A1N (.DIODE(_295_));
 scs8hd_diode_2 ANTENNA__607__A1 (.DIODE(_295_));
 scs8hd_diode_2 ANTENNA__608__A2N (.DIODE(_296_));
 scs8hd_diode_2 ANTENNA__607__A2 (.DIODE(_296_));
 scs8hd_diode_2 ANTENNA__626__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__619__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__612__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__605__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__338__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__331__A (.DIODE(_297_));
 scs8hd_diode_2 ANTENNA__606__A (.DIODE(_298_));
 scs8hd_diode_2 ANTENNA__609__A (.DIODE(_299_));
 scs8hd_diode_2 ANTENNA__608__B1 (.DIODE(_299_));
 scs8hd_diode_2 ANTENNA__609__B (.DIODE(_300_));
 scs8hd_diode_2 ANTENNA__608__B2 (.DIODE(_300_));
 scs8hd_diode_2 ANTENNA__615__A1N (.DIODE(_301_));
 scs8hd_diode_2 ANTENNA__614__A1 (.DIODE(_301_));
 scs8hd_diode_2 ANTENNA__615__A2N (.DIODE(_302_));
 scs8hd_diode_2 ANTENNA__614__A2 (.DIODE(_302_));
 scs8hd_diode_2 ANTENNA__613__A (.DIODE(_303_));
 scs8hd_diode_2 ANTENNA__616__A (.DIODE(_304_));
 scs8hd_diode_2 ANTENNA__615__B1 (.DIODE(_304_));
 scs8hd_diode_2 ANTENNA__616__B (.DIODE(_305_));
 scs8hd_diode_2 ANTENNA__615__B2 (.DIODE(_305_));
 scs8hd_diode_2 ANTENNA__622__A1N (.DIODE(_306_));
 scs8hd_diode_2 ANTENNA__621__A1 (.DIODE(_306_));
 scs8hd_diode_2 ANTENNA__622__A2N (.DIODE(_307_));
 scs8hd_diode_2 ANTENNA__621__A2 (.DIODE(_307_));
 scs8hd_diode_2 ANTENNA__620__A (.DIODE(_308_));
 scs8hd_diode_2 ANTENNA__623__A (.DIODE(_309_));
 scs8hd_diode_2 ANTENNA__622__B1 (.DIODE(_309_));
 scs8hd_diode_2 ANTENNA__623__B (.DIODE(_310_));
 scs8hd_diode_2 ANTENNA__622__B2 (.DIODE(_310_));
 scs8hd_diode_2 ANTENNA__629__A1N (.DIODE(_311_));
 scs8hd_diode_2 ANTENNA__628__A1 (.DIODE(_311_));
 scs8hd_diode_2 ANTENNA__629__A2N (.DIODE(_312_));
 scs8hd_diode_2 ANTENNA__628__A2 (.DIODE(_312_));
 scs8hd_diode_2 ANTENNA__627__A (.DIODE(_313_));
 scs8hd_diode_2 ANTENNA__630__A (.DIODE(_314_));
 scs8hd_diode_2 ANTENNA__629__B1 (.DIODE(_314_));
 scs8hd_diode_2 ANTENNA__630__B (.DIODE(_315_));
 scs8hd_diode_2 ANTENNA__629__B2 (.DIODE(_315_));
 scs8hd_diode_2 ANTENNA__334__A1N (.DIODE(_316_));
 scs8hd_diode_2 ANTENNA__333__A1 (.DIODE(_316_));
 scs8hd_diode_2 ANTENNA__334__A2N (.DIODE(_317_));
 scs8hd_diode_2 ANTENNA__333__A2 (.DIODE(_317_));
 scs8hd_diode_2 ANTENNA__332__A (.DIODE(_318_));
 scs8hd_diode_2 ANTENNA__335__A (.DIODE(_319_));
 scs8hd_diode_2 ANTENNA__334__B1 (.DIODE(_319_));
 scs8hd_diode_2 ANTENNA__335__B (.DIODE(_320_));
 scs8hd_diode_2 ANTENNA__334__B2 (.DIODE(_320_));
 scs8hd_diode_2 ANTENNA__341__A1N (.DIODE(_321_));
 scs8hd_diode_2 ANTENNA__340__A1 (.DIODE(_321_));
 scs8hd_diode_2 ANTENNA__341__A2N (.DIODE(_322_));
 scs8hd_diode_2 ANTENNA__340__A2 (.DIODE(_322_));
 scs8hd_diode_2 ANTENNA__339__A (.DIODE(_323_));
 scs8hd_diode_2 ANTENNA__342__A (.DIODE(_324_));
 scs8hd_diode_2 ANTENNA__341__B1 (.DIODE(_324_));
 scs8hd_diode_2 ANTENNA__342__B (.DIODE(_325_));
 scs8hd_diode_2 ANTENNA__341__B2 (.DIODE(_325_));
 scs8hd_diode_2 ANTENNA__348__A1N (.DIODE(_326_));
 scs8hd_diode_2 ANTENNA__347__A1 (.DIODE(_326_));
 scs8hd_diode_2 ANTENNA__348__A2N (.DIODE(_327_));
 scs8hd_diode_2 ANTENNA__347__A2 (.DIODE(_327_));
 scs8hd_diode_2 ANTENNA__346__A (.DIODE(_328_));
 scs8hd_diode_2 ANTENNA__349__A (.DIODE(_329_));
 scs8hd_diode_2 ANTENNA__348__B1 (.DIODE(_329_));
 scs8hd_diode_2 ANTENNA__349__B (.DIODE(_330_));
 scs8hd_diode_2 ANTENNA__348__B2 (.DIODE(_330_));
 scs8hd_diode_2 ANTENNA__648__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__647__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__646__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__645__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__644__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__643__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__642__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__641__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__640__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__639__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__638__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__637__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__636__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__635__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__634__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__633__CLK (.DIODE(clk_0_0));
 scs8hd_diode_2 ANTENNA__664__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__663__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__662__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__661__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__660__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__659__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__658__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__657__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__656__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__655__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__654__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__653__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__652__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__651__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__650__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__649__CLK (.DIODE(clk_0_16));
 scs8hd_diode_2 ANTENNA__680__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__679__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__678__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__677__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__676__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__675__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__674__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__673__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__672__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__671__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__670__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__669__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__668__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__667__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__666__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__665__CLK (.DIODE(clk_0_32));
 scs8hd_diode_2 ANTENNA__696__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__695__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__694__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__693__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__692__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__691__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__690__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__689__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__688__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__687__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__686__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__685__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__684__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__683__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__682__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__681__CLK (.DIODE(clk_0_48));
 scs8hd_diode_2 ANTENNA__CTS_buf_1_48_A (.DIODE(clk_1_0));
 scs8hd_diode_2 ANTENNA__CTS_buf_1_32_A (.DIODE(clk_1_0));
 scs8hd_diode_2 ANTENNA__CTS_buf_1_16_A (.DIODE(clk_1_0));
 scs8hd_diode_2 ANTENNA__CTS_buf_1_0_A (.DIODE(clk_1_0));
 scs8hd_diode_2 ANTENNA__634__D (.DIODE(\csa0.hsum2 ));
 scs8hd_diode_2 ANTENNA__432__B1 (.DIODE(\csa0.sc ));
 scs8hd_diode_2 ANTENNA__426__A (.DIODE(\csa0.sc ));
 scs8hd_diode_2 ANTENNA__432__B2 (.DIODE(\csa0.y ));
 scs8hd_diode_2 ANTENNA__427__A (.DIODE(\csa0.y ));
 scs8hd_diode_2 ANTENNA__499__B2 (.DIODE(\pp[10] ));
 scs8hd_diode_2 ANTENNA__496__A (.DIODE(\pp[10] ));
 scs8hd_diode_2 ANTENNA__506__B2 (.DIODE(\pp[11] ));
 scs8hd_diode_2 ANTENNA__503__A (.DIODE(\pp[11] ));
 scs8hd_diode_2 ANTENNA__513__B2 (.DIODE(\pp[12] ));
 scs8hd_diode_2 ANTENNA__510__A (.DIODE(\pp[12] ));
 scs8hd_diode_2 ANTENNA__521__B2 (.DIODE(\pp[13] ));
 scs8hd_diode_2 ANTENNA__517__A (.DIODE(\pp[13] ));
 scs8hd_diode_2 ANTENNA__528__B2 (.DIODE(\pp[14] ));
 scs8hd_diode_2 ANTENNA__525__A (.DIODE(\pp[14] ));
 scs8hd_diode_2 ANTENNA__535__B2 (.DIODE(\pp[15] ));
 scs8hd_diode_2 ANTENNA__532__A (.DIODE(\pp[15] ));
 scs8hd_diode_2 ANTENNA__542__B2 (.DIODE(\pp[16] ));
 scs8hd_diode_2 ANTENNA__539__A (.DIODE(\pp[16] ));
 scs8hd_diode_2 ANTENNA__549__B2 (.DIODE(\pp[17] ));
 scs8hd_diode_2 ANTENNA__546__A (.DIODE(\pp[17] ));
 scs8hd_diode_2 ANTENNA__556__B2 (.DIODE(\pp[18] ));
 scs8hd_diode_2 ANTENNA__553__A (.DIODE(\pp[18] ));
 scs8hd_diode_2 ANTENNA__564__B2 (.DIODE(\pp[19] ));
 scs8hd_diode_2 ANTENNA__560__A (.DIODE(\pp[19] ));
 scs8hd_diode_2 ANTENNA__571__B2 (.DIODE(\pp[20] ));
 scs8hd_diode_2 ANTENNA__568__A (.DIODE(\pp[20] ));
 scs8hd_diode_2 ANTENNA__578__B2 (.DIODE(\pp[21] ));
 scs8hd_diode_2 ANTENNA__575__A (.DIODE(\pp[21] ));
 scs8hd_diode_2 ANTENNA__585__B2 (.DIODE(\pp[22] ));
 scs8hd_diode_2 ANTENNA__582__A (.DIODE(\pp[22] ));
 scs8hd_diode_2 ANTENNA__592__B2 (.DIODE(\pp[23] ));
 scs8hd_diode_2 ANTENNA__589__A (.DIODE(\pp[23] ));
 scs8hd_diode_2 ANTENNA__599__B2 (.DIODE(\pp[24] ));
 scs8hd_diode_2 ANTENNA__596__A (.DIODE(\pp[24] ));
 scs8hd_diode_2 ANTENNA__607__B2 (.DIODE(\pp[25] ));
 scs8hd_diode_2 ANTENNA__603__A (.DIODE(\pp[25] ));
 scs8hd_diode_2 ANTENNA__614__B2 (.DIODE(\pp[26] ));
 scs8hd_diode_2 ANTENNA__611__A (.DIODE(\pp[26] ));
 scs8hd_diode_2 ANTENNA__621__B2 (.DIODE(\pp[27] ));
 scs8hd_diode_2 ANTENNA__618__A (.DIODE(\pp[27] ));
 scs8hd_diode_2 ANTENNA__628__B2 (.DIODE(\pp[28] ));
 scs8hd_diode_2 ANTENNA__625__A (.DIODE(\pp[28] ));
 scs8hd_diode_2 ANTENNA__632__A (.DIODE(\pp[29] ));
 scs8hd_diode_2 ANTENNA__333__B2 (.DIODE(\pp[29] ));
 scs8hd_diode_2 ANTENNA__442__B2 (.DIODE(\pp[2] ));
 scs8hd_diode_2 ANTENNA__439__A (.DIODE(\pp[2] ));
 scs8hd_diode_2 ANTENNA__340__B2 (.DIODE(\pp[30] ));
 scs8hd_diode_2 ANTENNA__337__A (.DIODE(\pp[30] ));
 scs8hd_diode_2 ANTENNA__449__B2 (.DIODE(\pp[3] ));
 scs8hd_diode_2 ANTENNA__446__A (.DIODE(\pp[3] ));
 scs8hd_diode_2 ANTENNA__456__B2 (.DIODE(\pp[4] ));
 scs8hd_diode_2 ANTENNA__453__A (.DIODE(\pp[4] ));
 scs8hd_diode_2 ANTENNA__463__B2 (.DIODE(\pp[5] ));
 scs8hd_diode_2 ANTENNA__460__A (.DIODE(\pp[5] ));
 scs8hd_diode_2 ANTENNA__470__B2 (.DIODE(\pp[6] ));
 scs8hd_diode_2 ANTENNA__467__A (.DIODE(\pp[6] ));
 scs8hd_diode_2 ANTENNA__478__B2 (.DIODE(\pp[7] ));
 scs8hd_diode_2 ANTENNA__474__A (.DIODE(\pp[7] ));
 scs8hd_diode_2 ANTENNA__485__B2 (.DIODE(\pp[8] ));
 scs8hd_diode_2 ANTENNA__482__A (.DIODE(\pp[8] ));
 scs8hd_diode_2 ANTENNA__492__B2 (.DIODE(\pp[9] ));
 scs8hd_diode_2 ANTENNA__489__A (.DIODE(\pp[9] ));
 scs8hd_diode_2 ANTENNA__347__B2 (.DIODE(\tcmp.s ));
 scs8hd_diode_2 ANTENNA__344__A (.DIODE(\tcmp.s ));
 scs8hd_diode_2 ANTENNA__437__A1 (.DIODE(\tcmp.z ));
 scs8hd_diode_2 ANTENNA__436__A (.DIODE(\tcmp.z ));
endmodule
