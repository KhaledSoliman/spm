* NGSPICE file created from spm.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_4 abstract view
.subckt scs8hd_clkbuf_4 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_xor2_4 abstract view
.subckt scs8hd_xor2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_o22a_4 abstract view
.subckt scs8hd_o22a_4 A1 A2 B1 B2 X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfrtp_4 abstract view
.subckt scs8hd_dfrtp_4 CLK D Q RESETB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_a2bb2o_4 abstract view
.subckt scs8hd_a2bb2o_4 A1N A2N B1 B2 X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and2_4 abstract view
.subckt scs8hd_and2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_clkbuf_16 abstract view
.subckt scs8hd_clkbuf_16 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_a21boi_4 abstract view
.subckt scs8hd_a21boi_4 A1 A2 B1N Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt spm clk p rst x[0] x[10] x[11] x[12] x[13] x[14] x[15] x[16] x[17] x[18] x[19]
+ x[1] x[20] x[21] x[22] x[23] x[24] x[25] x[26] x[27] x[28] x[29] x[2] x[30] x[31]
+ x[3] x[4] x[5] x[6] x[7] x[8] x[9] y VDD VSS
XANTENNA__666__D _544_/X VSS VDD scs8hd_diode_2
XANTENNA__586__B2 _587_/B VSS VDD scs8hd_diode_2
XFILLER_22_100 VSS VDD scs8hd_decap_4
X_CTS_buf_1_16 _CTS_root/X _651_/CLK VSS VDD scs8hd_clkbuf_4
X_501_ _498_/X _501_/B _501_/X VSS VDD scs8hd_xor2_4
XANTENNA__682__RESETB _368_/X VSS VDD scs8hd_diode_2
XFILLER_26_41 VSS VDD scs8hd_decap_3
X_432_ _426_/Y _427_/Y _633_/Q _638_/Q _434_/B VSS VDD scs8hd_o22a_4
XFILLER_13_100 VDD VSS scs8hd_fill_2
XFILLER_42_40 VSS VDD scs8hd_fill_1
X_363_ _363_/A _363_/X VSS VDD scs8hd_buf_1
XFILLER_13_188 VDD VSS scs8hd_fill_2
XFILLER_3_56 VSS VDD scs8hd_fill_1
XFILLER_3_89 VSS VDD scs8hd_decap_4
XFILLER_8_170 VDD VSS scs8hd_fill_2
XANTENNA__633__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_6_118 VSS VDD scs8hd_decap_4
XFILLER_12_32 VDD VSS scs8hd_fill_2
XFILLER_12_76 VSS VDD scs8hd_decap_4
XFILLER_37_62 VSS VDD scs8hd_decap_3
XFILLER_37_51 VDD VSS scs8hd_fill_2
XFILLER_33_228 VDD VSS scs8hd_fill_2
X_346_ _345_/X _346_/X VSS VDD scs8hd_buf_1
X_415_ _410_/A _415_/X VSS VDD scs8hd_buf_1
XANTENNA__656__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_5_162 VDD VSS scs8hd_fill_2
XANTENNA__486__B1 _484_/X VSS VDD scs8hd_diode_2
XFILLER_5_184 VDD VSS scs8hd_fill_2
XFILLER_24_206 VDD VSS scs8hd_fill_2
XFILLER_32_250 VSS VDD scs8hd_decap_3
XFILLER_15_206 VDD VSS scs8hd_fill_2
XFILLER_15_217 VDD VSS scs8hd_fill_2
XFILLER_15_228 VDD VSS scs8hd_fill_2
XANTENNA__679__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_2_165 VSS VDD scs8hd_decap_6
XFILLER_2_154 VDD VSS scs8hd_fill_2
XFILLER_0_24 VSS VDD scs8hd_decap_3
XFILLER_9_99 VSS VDD scs8hd_decap_4
XFILLER_14_250 VSS VDD scs8hd_decap_3
XFILLER_21_209 VSS VDD scs8hd_decap_4
XANTENNA__471__A2N _467_/Y VSS VDD scs8hd_diode_2
XANTENNA__674__D _674_/D VSS VDD scs8hd_diode_2
X_680_ _667_/CLK _680_/D _582_/A _370_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__622__B1 _623_/A VSS VDD scs8hd_diode_2
XFILLER_18_20 VDD VSS scs8hd_fill_2
XFILLER_11_220 VDD VSS scs8hd_fill_2
XFILLER_38_106 VDD VSS scs8hd_fill_2
XANTENNA__402__A _402_/A VSS VDD scs8hd_diode_2
XANTENNA__669__D _669_/D VSS VDD scs8hd_diode_2
XFILLER_37_172 VSS VDD scs8hd_decap_3
XFILLER_37_161 VDD VSS scs8hd_fill_2
XFILLER_4_205 VSS VDD scs8hd_fill_1
XFILLER_20_32 VSS VDD scs8hd_decap_3
XFILLER_29_85 VDD VSS scs8hd_fill_2
XFILLER_29_52 VDD VSS scs8hd_fill_2
XFILLER_20_87 VSS VDD scs8hd_fill_1
X_663_ _651_/CLK _536_/X _663_/Q _391_/X VSS VDD scs8hd_dfrtp_4
X_594_ _594_/A _592_/X _680_/D VSS VDD scs8hd_xor2_4
XFILLER_28_183 VDD VSS scs8hd_fill_2
XFILLER_6_23 VDD VSS scs8hd_fill_2
XANTENNA__677__RESETB _375_/X VSS VDD scs8hd_diode_2
XANTENNA__565__A1N _559_/Y VSS VDD scs8hd_diode_2
XFILLER_13_3 VDD VSS scs8hd_fill_2
XFILLER_19_172 VSS VDD scs8hd_decap_3
XFILLER_25_153 VDD VSS scs8hd_fill_2
XFILLER_31_53 VDD VSS scs8hd_fill_2
XFILLER_31_31 VSS VDD scs8hd_decap_4
XFILLER_15_87 VDD VSS scs8hd_fill_2
XFILLER_31_123 VSS VDD scs8hd_decap_4
XANTENNA__347__A2 _344_/Y VSS VDD scs8hd_diode_2
X_646_ _648_/CLK _472_/X _460_/A _411_/X VSS VDD scs8hd_dfrtp_4
X_577_ _577_/A _580_/A VSS VDD scs8hd_buf_1
XPHY_170 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_192 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_181 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_39_245 VSS VDD scs8hd_decap_8
XANTENNA__682__D _601_/X VSS VDD scs8hd_diode_2
XFILLER_22_145 VSS VDD scs8hd_decap_4
XFILLER_7_8 VDD VSS scs8hd_fill_2
X_500_ _495_/Y _496_/Y _498_/X _501_/B _653_/D VSS VDD scs8hd_a2bb2o_4
XFILLER_26_64 VDD VSS scs8hd_fill_2
X_431_ _431_/A _434_/A VSS VDD scs8hd_buf_1
X_362_ _363_/A _362_/X VSS VDD scs8hd_buf_1
XFILLER_13_112 VDD VSS scs8hd_fill_2
XFILLER_13_123 VDD VSS scs8hd_fill_2
XFILLER_42_85 VSS VDD scs8hd_decap_8
XFILLER_42_63 VSS VDD scs8hd_decap_12
XFILLER_42_52 VSS VDD scs8hd_decap_8
XFILLER_13_178 VSS VDD scs8hd_decap_4
XANTENNA__410__A _410_/A VSS VDD scs8hd_diode_2
XFILLER_36_215 VDD VSS scs8hd_fill_2
X_629_ _624_/Y _625_/Y _627_/X _630_/B _629_/X VSS VDD scs8hd_a2bb2o_4
XANTENNA__677__D _586_/X VSS VDD scs8hd_diode_2
XFILLER_42_218 VSS VDD scs8hd_decap_12
XFILLER_10_159 VSS VDD scs8hd_decap_4
XFILLER_37_41 VDD VSS scs8hd_fill_2
XFILLER_18_215 VSS VDD scs8hd_decap_4
XFILLER_41_240 VSS VDD scs8hd_decap_4
X_345_ _518_/A x[30] _345_/X VSS VDD scs8hd_and2_4
X_414_ _410_/A _414_/X VSS VDD scs8hd_buf_1
XANTENNA__405__A _405_/A VSS VDD scs8hd_diode_2
XFILLER_5_141 VSS VDD scs8hd_decap_4
XANTENNA__486__B2 _485_/X VSS VDD scs8hd_diode_2
XFILLER_24_229 VSS VDD scs8hd_decap_4
XFILLER_23_54 VDD VSS scs8hd_fill_2
XFILLER_23_10 VDD VSS scs8hd_fill_2
XFILLER_23_87 VDD VSS scs8hd_fill_2
XFILLER_23_76 VSS VDD scs8hd_decap_4
XFILLER_2_122 VSS VDD scs8hd_decap_3
XFILLER_9_23 VDD VSS scs8hd_fill_2
XFILLER_9_67 VDD VSS scs8hd_fill_2
XANTENNA__471__A1N _466_/Y VSS VDD scs8hd_diode_2
XANTENNA__690__D _630_/X VSS VDD scs8hd_diode_2
XANTENNA__622__B2 _623_/B VSS VDD scs8hd_diode_2
XANTENNA__646__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_18_32 VSS VDD scs8hd_decap_8
XFILLER_34_86 VDD VSS scs8hd_fill_2
XFILLER_34_75 VSS VDD scs8hd_decap_4
XFILLER_7_236 VDD VSS scs8hd_fill_2
XFILLER_11_243 VSS VDD scs8hd_fill_1
XANTENNA__673__RESETB _379_/X VSS VDD scs8hd_diode_2
XFILLER_37_184 VSS VDD scs8hd_decap_4
XANTENNA__669__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_1_90 VDD VSS scs8hd_fill_2
XANTENNA__685__D _685_/D VSS VDD scs8hd_diode_2
XANTENNA__503__A _658_/Q VSS VDD scs8hd_diode_2
XFILLER_28_140 VSS VDD scs8hd_decap_4
X_662_ _651_/CLK _662_/D _662_/Q _392_/X VSS VDD scs8hd_dfrtp_4
X_593_ _588_/Y _589_/Y _594_/A _592_/X _593_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_28_195 VDD VSS scs8hd_fill_2
XFILLER_28_151 VDD VSS scs8hd_fill_2
XFILLER_6_57 VDD VSS scs8hd_fill_2
XFILLER_6_79 VDD VSS scs8hd_fill_2
XANTENNA__413__A _410_/A VSS VDD scs8hd_diode_2
XFILLER_19_140 VDD VSS scs8hd_fill_2
XFILLER_19_184 VDD VSS scs8hd_fill_2
XFILLER_34_154 VSS VDD scs8hd_decap_8
XANTENNA__522__B1 _520_/X VSS VDD scs8hd_diode_2
XFILLER_25_132 VSS VDD scs8hd_decap_8
XFILLER_25_121 VSS VDD scs8hd_fill_1
XFILLER_15_55 VDD VSS scs8hd_fill_2
XANTENNA__334__A2N _632_/Y VSS VDD scs8hd_diode_2
XANTENNA__513__B1 _657_/Q VSS VDD scs8hd_diode_2
X_645_ _648_/CLK _471_/X _645_/Q _412_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__408__A _405_/A VSS VDD scs8hd_diode_2
XPHY_193 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_182 VSS VDD scs8hd_tapvpwrvgnd_1
X_576_ _597_/A x[20] _577_/A VSS VDD scs8hd_and2_4
XFILLER_16_154 VDD VSS scs8hd_fill_2
XPHY_160 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_171 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_39_235 VDD VSS scs8hd_fill_2
XFILLER_30_190 VSS VDD scs8hd_decap_4
XFILLER_22_179 VSS VDD scs8hd_decap_4
XFILLER_22_135 VSS VDD scs8hd_decap_6
XFILLER_26_32 VSS VDD scs8hd_decap_3
XFILLER_26_21 VDD VSS scs8hd_fill_2
XFILLER_26_98 VSS VDD scs8hd_decap_6
X_430_ _461_/A x[0] _431_/A VSS VDD scs8hd_and2_4
XFILLER_9_139 VDD VSS scs8hd_fill_2
X_361_ _363_/A _361_/X VSS VDD scs8hd_buf_1
XFILLER_42_75 VSS VDD scs8hd_decap_3
XFILLER_36_205 VSS VDD scs8hd_decap_4
X_628_ _624_/Y _625_/Y _624_/A _625_/A _630_/B VSS VDD scs8hd_o22a_4
X_559_ _671_/Q _559_/Y VSS VDD scs8hd_inv_8
XANTENNA__601__A _598_/X VSS VDD scs8hd_diode_2
XFILLER_8_194 VDD VSS scs8hd_fill_2
XANTENNA__693__D _341_/X VSS VDD scs8hd_diode_2
XFILLER_10_127 VSS VDD scs8hd_decap_12
XFILLER_12_12 VSS VDD scs8hd_decap_4
XFILLER_12_23 VDD VSS scs8hd_fill_2
X_CTS_buf_1_0 _CTS_root/X _648_/CLK VSS VDD scs8hd_clkbuf_4
XANTENNA__511__A _476_/A VSS VDD scs8hd_diode_2
XANTENNA__522__A2N _517_/Y VSS VDD scs8hd_diode_2
XFILLER_37_97 VDD VSS scs8hd_fill_2
X_413_ _410_/A _413_/X VSS VDD scs8hd_buf_1
X_344_ _344_/A _344_/Y VSS VDD scs8hd_inv_8
XANTENNA__421__A _417_/A VSS VDD scs8hd_diode_2
XANTENNA__668__RESETB _385_/X VSS VDD scs8hd_diode_2
XANTENNA__331__A _605_/A VSS VDD scs8hd_diode_2
XANTENNA__688__D _688_/D VSS VDD scs8hd_diode_2
XFILLER_23_66 VSS VDD scs8hd_decap_3
XFILLER_3_3 VSS VDD scs8hd_decap_12
XFILLER_2_145 VSS VDD scs8hd_decap_4
XFILLER_0_37 VDD VSS scs8hd_fill_2
XFILLER_9_35 VDD VSS scs8hd_fill_2
XANTENNA__416__A _373_/A VSS VDD scs8hd_diode_2
XFILLER_9_57 VSS VDD scs8hd_decap_4
XFILLER_36_3 VDD VSS scs8hd_fill_2
XFILLER_18_44 VDD VSS scs8hd_fill_2
XFILLER_34_32 VDD VSS scs8hd_fill_2
XFILLER_34_21 VDD VSS scs8hd_fill_2
XFILLER_18_66 VSS VDD scs8hd_fill_1
XFILLER_18_99 VDD VSS scs8hd_fill_2
XFILLER_7_215 VSS VDD scs8hd_fill_1
XFILLER_11_233 VDD VSS scs8hd_fill_2
XFILLER_37_130 VDD VSS scs8hd_fill_2
XFILLER_29_10 VDD VSS scs8hd_fill_2
XFILLER_4_229 VDD VSS scs8hd_fill_2
X_592_ _588_/Y _589_/Y _679_/Q _682_/Q _592_/X VSS VDD scs8hd_o22a_4
X_661_ _651_/CLK _661_/D _661_/Q _393_/X VSS VDD scs8hd_dfrtp_4
XFILLER_29_76 VDD VSS scs8hd_fill_2
XFILLER_28_174 VDD VSS scs8hd_fill_2
XFILLER_34_188 VDD VSS scs8hd_fill_2
XANTENNA__604__A y VSS VDD scs8hd_diode_2
XANTENNA__636__CLK _648_/CLK VSS VDD scs8hd_diode_2
XANTENNA__522__B2 _521_/X VSS VDD scs8hd_diode_2
XANTENNA__696__D _349_/X VSS VDD scs8hd_diode_2
XFILLER_40_158 VSS VDD scs8hd_fill_1
XFILLER_40_147 VDD VSS scs8hd_fill_2
XFILLER_40_125 VDD VSS scs8hd_fill_2
XFILLER_25_144 VDD VSS scs8hd_fill_2
XFILLER_25_100 VDD VSS scs8hd_fill_2
XANTENNA__334__A1N _631_/Y VSS VDD scs8hd_diode_2
XFILLER_31_88 VSS VDD scs8hd_decap_4
XFILLER_31_77 VSS VDD scs8hd_decap_4
XANTENNA__513__A1 _509_/Y VSS VDD scs8hd_diode_2
XANTENNA__629__A2N _625_/Y VSS VDD scs8hd_diode_2
XANTENNA__513__B2 _660_/Q VSS VDD scs8hd_diode_2
X_575_ _678_/Q _575_/Y VSS VDD scs8hd_inv_8
X_644_ _648_/CLK _465_/X _644_/Q _413_/X VSS VDD scs8hd_dfrtp_4
XFILLER_31_114 VSS VDD scs8hd_decap_4
XPHY_194 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_183 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__659__CLK _651_/CLK VSS VDD scs8hd_diode_2
XANTENNA__424__A _366_/A VSS VDD scs8hd_diode_2
XPHY_150 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_161 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_172 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__509__A _657_/Q VSS VDD scs8hd_diode_2
XFILLER_42_32 VSS VDD scs8hd_decap_8
X_360_ _363_/A _360_/X VSS VDD scs8hd_buf_1
XFILLER_42_98 VSS VDD scs8hd_decap_6
XFILLER_3_59 VDD VSS scs8hd_fill_2
XFILLER_3_48 VDD VSS scs8hd_fill_2
XFILLER_3_15 VSS VDD scs8hd_fill_1
XFILLER_36_239 VDD VSS scs8hd_fill_2
X_558_ _558_/A _558_/B _670_/D VSS VDD scs8hd_xor2_4
XANTENNA__419__A _417_/A VSS VDD scs8hd_diode_2
X_627_ _626_/X _627_/X VSS VDD scs8hd_buf_1
X_489_ _489_/A _489_/Y VSS VDD scs8hd_inv_8
XFILLER_8_151 VDD VSS scs8hd_fill_2
XANTENNA__601__B _601_/B VSS VDD scs8hd_diode_2
XANTENNA__664__RESETB _390_/X VSS VDD scs8hd_diode_2
XFILLER_27_239 VSS VDD scs8hd_decap_4
XFILLER_10_139 VDD VSS scs8hd_fill_2
XFILLER_12_46 VSS VDD scs8hd_decap_4
XFILLER_12_57 VDD VSS scs8hd_fill_2
XANTENNA__511__B x[11] VSS VDD scs8hd_diode_2
XFILLER_18_206 VSS VDD scs8hd_decap_4
XANTENNA__522__A1N _516_/Y VSS VDD scs8hd_diode_2
X_412_ _410_/A _412_/X VSS VDD scs8hd_buf_1
XFILLER_5_121 VSS VDD scs8hd_fill_1
X_343_ _343_/A _343_/Y VSS VDD scs8hd_inv_8
XFILLER_5_154 VDD VSS scs8hd_fill_2
XFILLER_5_176 VSS VDD scs8hd_decap_3
XFILLER_32_242 VSS VDD scs8hd_decap_8
XFILLER_32_220 VDD VSS scs8hd_fill_2
XANTENNA__612__A _605_/A VSS VDD scs8hd_diode_2
XANTENNA__331__B x[28] VSS VDD scs8hd_diode_2
XFILLER_23_242 VDD VSS scs8hd_fill_2
XFILLER_0_49 VSS VDD scs8hd_decap_12
XFILLER_14_220 VDD VSS scs8hd_fill_2
XFILLER_14_242 VSS VDD scs8hd_decap_8
XFILLER_29_3 VSS VDD scs8hd_decap_4
XFILLER_20_201 VDD VSS scs8hd_fill_2
XFILLER_20_212 VDD VSS scs8hd_fill_2
XANTENNA__342__A _339_/X VSS VDD scs8hd_diode_2
XANTENNA__607__B1 _683_/Q VSS VDD scs8hd_diode_2
XFILLER_18_12 VDD VSS scs8hd_fill_2
XANTENNA__517__A _662_/Q VSS VDD scs8hd_diode_2
XFILLER_18_78 VSS VDD scs8hd_decap_12
XANTENNA__692__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_7_249 VSS VDD scs8hd_decap_4
XFILLER_11_245 VSS VDD scs8hd_decap_8
XANTENNA__427__A _638_/Q VSS VDD scs8hd_diode_2
XFILLER_37_120 VDD VSS scs8hd_fill_2
XANTENNA__337__A _337_/A VSS VDD scs8hd_diode_2
XFILLER_4_208 VDD VSS scs8hd_fill_2
XFILLER_20_24 VDD VSS scs8hd_fill_2
XFILLER_29_44 VDD VSS scs8hd_fill_2
XFILLER_20_57 VSS VDD scs8hd_decap_4
X_591_ _590_/X _594_/A VSS VDD scs8hd_buf_1
XFILLER_28_131 VSS VDD scs8hd_decap_6
X_660_ _651_/CLK _660_/D _660_/Q _394_/X VSS VDD scs8hd_dfrtp_4
XFILLER_3_230 VDD VSS scs8hd_fill_2
XFILLER_10_90 VDD VSS scs8hd_fill_2
XFILLER_20_7 VSS VDD scs8hd_decap_4
XFILLER_19_120 VDD VSS scs8hd_fill_2
XFILLER_19_131 VSS VDD scs8hd_decap_6
XFILLER_34_145 VDD VSS scs8hd_fill_2
XFILLER_34_134 VSS VDD scs8hd_decap_8
XFILLER_34_123 VDD VSS scs8hd_fill_2
XFILLER_19_164 VDD VSS scs8hd_fill_2
XANTENNA__620__A _620_/A VSS VDD scs8hd_diode_2
XFILLER_25_123 VDD VSS scs8hd_fill_2
XFILLER_25_178 VSS VDD scs8hd_fill_1
XANTENNA__513__A2 _510_/Y VSS VDD scs8hd_diode_2
XANTENNA__629__A1N _624_/Y VSS VDD scs8hd_diode_2
XANTENNA__659__RESETB _396_/X VSS VDD scs8hd_diode_2
XANTENNA__530__A _527_/X VSS VDD scs8hd_diode_2
XFILLER_0_222 VDD VSS scs8hd_fill_2
X_574_ _574_/A _574_/Y VSS VDD scs8hd_inv_8
X_643_ _648_/CLK _643_/D _643_/Q _414_/X VSS VDD scs8hd_dfrtp_4
XPHY_195 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_184 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_140 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_151 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_162 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_173 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__440__A _461_/A VSS VDD scs8hd_diode_2
XFILLER_11_3 VDD VSS scs8hd_fill_2
XFILLER_30_170 VSS VDD scs8hd_decap_3
XFILLER_7_91 VSS VDD scs8hd_decap_4
XANTENNA__660__RESETB _394_/X VSS VDD scs8hd_diode_2
XANTENNA__350__A _366_/A VSS VDD scs8hd_diode_2
XFILLER_13_104 VDD VSS scs8hd_fill_2
XANTENNA__525__A _664_/Q VSS VDD scs8hd_diode_2
XFILLER_13_148 VDD VSS scs8hd_fill_2
XFILLER_21_170 VSS VDD scs8hd_decap_4
XFILLER_21_181 VDD VSS scs8hd_fill_2
X_488_ _488_/A _488_/Y VSS VDD scs8hd_inv_8
X_557_ _552_/Y _553_/Y _558_/A _558_/B _669_/D VSS VDD scs8hd_a2bb2o_4
X_626_ _605_/A x[27] _626_/X VSS VDD scs8hd_and2_4
XANTENNA__435__A _518_/A VSS VDD scs8hd_diode_2
XFILLER_8_174 VDD VSS scs8hd_fill_2
XFILLER_35_240 VSS VDD scs8hd_decap_4
XFILLER_10_118 VSS VDD scs8hd_decap_3
XANTENNA__345__A _518_/A VSS VDD scs8hd_diode_2
XFILLER_12_36 VDD VSS scs8hd_fill_2
XFILLER_37_55 VDD VSS scs8hd_fill_2
XANTENNA__649__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_41_221 VSS VDD scs8hd_decap_4
X_342_ _339_/X _340_/X _694_/D VSS VDD scs8hd_xor2_4
X_411_ _410_/A _411_/X VSS VDD scs8hd_buf_1
XFILLER_5_133 VDD VSS scs8hd_fill_2
XFILLER_38_8 VSS VDD scs8hd_decap_3
XANTENNA__340__B1 _693_/Q VSS VDD scs8hd_diode_2
XFILLER_5_166 VSS VDD scs8hd_decap_3
X_609_ _609_/A _609_/B _684_/D VSS VDD scs8hd_xor2_4
XFILLER_17_240 VSS VDD scs8hd_decap_4
XFILLER_32_232 VSS VDD scs8hd_fill_1
XANTENNA__612__B x[25] VSS VDD scs8hd_diode_2
XFILLER_4_70 VDD VSS scs8hd_fill_2
XFILLER_23_46 VDD VSS scs8hd_fill_2
XFILLER_23_35 VSS VDD scs8hd_decap_3
XANTENNA__464__A2N _460_/Y VSS VDD scs8hd_diode_2
XFILLER_1_191 VDD VSS scs8hd_fill_2
XANTENNA__623__A _623_/A VSS VDD scs8hd_diode_2
XANTENNA__342__B _340_/X VSS VDD scs8hd_diode_2
XANTENNA__607__B2 _603_/A VSS VDD scs8hd_diode_2
XANTENNA__607__A1 _602_/Y VSS VDD scs8hd_diode_2
XFILLER_18_24 VSS VDD scs8hd_decap_3
XFILLER_34_45 VSS VDD scs8hd_fill_1
XFILLER_11_213 VSS VDD scs8hd_fill_1
XANTENNA__533__A _547_/A VSS VDD scs8hd_diode_2
XANTENNA__543__B1 _544_/A VSS VDD scs8hd_diode_2
XFILLER_41_3 VSS VDD scs8hd_decap_12
XANTENNA__618__A _690_/Q VSS VDD scs8hd_diode_2
XANTENNA__353__A _357_/A VSS VDD scs8hd_diode_2
XFILLER_29_67 VDD VSS scs8hd_fill_2
XFILLER_29_56 VSS VDD scs8hd_decap_4
X_590_ _597_/A x[22] _590_/X VSS VDD scs8hd_and2_4
XFILLER_29_89 VDD VSS scs8hd_fill_2
XFILLER_28_187 VSS VDD scs8hd_decap_4
XFILLER_28_154 VDD VSS scs8hd_fill_2
XFILLER_28_110 VSS VDD scs8hd_decap_3
XANTENNA__655__RESETB _400_/X VSS VDD scs8hd_diode_2
XFILLER_6_27 VSS VDD scs8hd_decap_4
XFILLER_13_7 VDD VSS scs8hd_fill_2
XFILLER_34_113 VSS VDD scs8hd_decap_3
XANTENNA__438__A _438_/A VSS VDD scs8hd_diode_2
XANTENNA__507__B1 _508_/A VSS VDD scs8hd_diode_2
XANTENNA__682__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_25_157 VDD VSS scs8hd_fill_2
XFILLER_25_113 VDD VSS scs8hd_fill_2
XFILLER_25_168 VDD VSS scs8hd_fill_2
XFILLER_15_47 VDD VSS scs8hd_fill_2
XFILLER_31_57 VSS VDD scs8hd_decap_4
XANTENNA__530__B _528_/X VSS VDD scs8hd_diode_2
XFILLER_0_245 VSS VDD scs8hd_decap_3
X_642_ _648_/CLK _458_/X _446_/A _415_/X VSS VDD scs8hd_dfrtp_4
XFILLER_31_149 VSS VDD scs8hd_decap_4
XPHY_130 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_141 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_152 VSS VDD scs8hd_tapvpwrvgnd_1
X_573_ _570_/X _573_/B _674_/D VSS VDD scs8hd_xor2_4
XPHY_196 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_185 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_163 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_174 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_39_216 VDD VSS scs8hd_fill_2
XANTENNA__440__B x[1] VSS VDD scs8hd_diode_2
XFILLER_39_227 VDD VSS scs8hd_fill_2
XANTENNA__631__A _691_/Q VSS VDD scs8hd_diode_2
XFILLER_26_68 VSS VDD scs8hd_decap_12
XFILLER_26_13 VDD VSS scs8hd_fill_2
XFILLER_13_116 VDD VSS scs8hd_fill_2
XFILLER_21_193 VDD VSS scs8hd_fill_2
XANTENNA__541__A _540_/X VSS VDD scs8hd_diode_2
X_625_ _625_/A _625_/Y VSS VDD scs8hd_inv_8
X_487_ _484_/X _485_/X _487_/X VSS VDD scs8hd_xor2_4
X_556_ _552_/Y _553_/Y _552_/A _553_/A _558_/B VSS VDD scs8hd_o22a_4
XFILLER_12_171 VSS VDD scs8hd_decap_4
XANTENNA__435__B x[31] VSS VDD scs8hd_diode_2
XFILLER_16_90 VDD VSS scs8hd_fill_2
XANTENNA__451__A _451_/A VSS VDD scs8hd_diode_2
XFILLER_12_182 VSS VDD scs8hd_decap_3
XANTENNA__626__A _605_/A VSS VDD scs8hd_diode_2
XANTENNA__345__B x[30] VSS VDD scs8hd_diode_2
XANTENNA__361__A _363_/A VSS VDD scs8hd_diode_2
XFILLER_37_67 VDD VSS scs8hd_fill_2
XFILLER_37_45 VSS VDD scs8hd_decap_3
XFILLER_37_34 VSS VDD scs8hd_decap_4
XFILLER_18_219 VSS VDD scs8hd_fill_1
X_341_ _336_/Y _337_/Y _339_/X _340_/X _341_/X VSS VDD scs8hd_a2bb2o_4
X_410_ _410_/A _410_/X VSS VDD scs8hd_buf_1
XFILLER_5_123 VDD VSS scs8hd_fill_2
XANTENNA__340__A1 _336_/Y VSS VDD scs8hd_diode_2
XANTENNA__340__B2 _337_/A VSS VDD scs8hd_diode_2
X_608_ _602_/Y _603_/Y _609_/A _609_/B _683_/D VSS VDD scs8hd_a2bb2o_4
XANTENNA__446__A _446_/A VSS VDD scs8hd_diode_2
XANTENNA__CTS_root_A clk VSS VDD scs8hd_diode_2
X_539_ _539_/A _539_/Y VSS VDD scs8hd_inv_8
XFILLER_4_93 VDD VSS scs8hd_fill_2
XANTENNA__356__A _357_/A VSS VDD scs8hd_diode_2
XFILLER_23_58 VSS VDD scs8hd_decap_3
XFILLER_0_29 VDD VSS scs8hd_fill_2
XFILLER_9_27 VSS VDD scs8hd_decap_4
XANTENNA__464__A1N _459_/Y VSS VDD scs8hd_diode_2
XFILLER_1_170 VDD VSS scs8hd_fill_2
XANTENNA__639__CLK _648_/CLK VSS VDD scs8hd_diode_2
XANTENNA__623__B _623_/B VSS VDD scs8hd_diode_2
XANTENNA__607__A2 _603_/Y VSS VDD scs8hd_diode_2
XFILLER_18_69 VDD VSS scs8hd_fill_2
XFILLER_34_79 VSS VDD scs8hd_fill_1
XFILLER_7_218 VDD VSS scs8hd_fill_2
XANTENNA__533__B x[14] VSS VDD scs8hd_diode_2
XANTENNA__543__B2 _544_/B VSS VDD scs8hd_diode_2
XANTENNA__651__RESETB _405_/X VSS VDD scs8hd_diode_2
XFILLER_1_3 VSS VDD scs8hd_decap_3
XFILLER_34_3 VDD VSS scs8hd_fill_2
XFILLER_37_177 VDD VSS scs8hd_fill_2
XFILLER_37_155 VSS VDD scs8hd_decap_4
XANTENNA__470__B1 _645_/Q VSS VDD scs8hd_diode_2
XFILLER_29_35 VDD VSS scs8hd_fill_2
XFILLER_28_199 VDD VSS scs8hd_fill_2
XFILLER_28_144 VSS VDD scs8hd_fill_1
XANTENNA__544__A _544_/A VSS VDD scs8hd_diode_2
XFILLER_19_177 VDD VSS scs8hd_fill_2
XANTENNA__454__A _461_/A VSS VDD scs8hd_diode_2
XANTENNA__507__B2 _508_/B VSS VDD scs8hd_diode_2
XANTENNA__443__B1 _441_/X VSS VDD scs8hd_diode_2
XFILLER_15_59 VDD VSS scs8hd_fill_2
XANTENNA__364__A _363_/A VSS VDD scs8hd_diode_2
XFILLER_0_213 VSS VDD scs8hd_decap_4
XANTENNA__539__A _539_/A VSS VDD scs8hd_diode_2
X_641_ _648_/CLK _457_/X _452_/A _417_/X VSS VDD scs8hd_dfrtp_4
X_572_ _567_/Y _568_/Y _570_/X _573_/B _572_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_16_103 VDD VSS scs8hd_fill_2
XFILLER_24_191 VSS VDD scs8hd_decap_4
XPHY_120 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_131 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_142 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_153 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_16_125 VSS VDD scs8hd_decap_8
XFILLER_16_147 VDD VSS scs8hd_fill_2
XFILLER_16_169 VSS VDD scs8hd_fill_1
XPHY_164 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_175 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_197 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_186 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_21_91 VDD VSS scs8hd_fill_2
XFILLER_39_239 VSS VDD scs8hd_decap_4
XFILLER_22_106 VDD VSS scs8hd_fill_2
XPHY_0 VSS VDD scs8hd_decap_3
XFILLER_30_194 VSS VDD scs8hd_fill_1
XFILLER_30_183 VSS VDD scs8hd_fill_1
XFILLER_7_82 VDD VSS scs8hd_fill_2
XANTENNA__359__A _366_/A VSS VDD scs8hd_diode_2
XFILLER_26_25 VDD VSS scs8hd_fill_2
XFILLER_21_150 VDD VSS scs8hd_fill_2
XFILLER_3_18 VDD VSS scs8hd_fill_2
XFILLER_36_209 VSS VDD scs8hd_fill_1
X_555_ _554_/X _558_/A VSS VDD scs8hd_buf_1
X_624_ _624_/A _624_/Y VSS VDD scs8hd_inv_8
X_486_ _481_/Y _482_/Y _484_/X _485_/X _486_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_8_143 VDD VSS scs8hd_fill_2
XFILLER_8_154 VDD VSS scs8hd_fill_2
XFILLER_32_90 VDD VSS scs8hd_fill_2
XANTENNA__672__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__451__B _449_/X VSS VDD scs8hd_diode_2
XFILLER_8_198 VSS VDD scs8hd_decap_4
XFILLER_27_209 VDD VSS scs8hd_fill_2
XFILLER_35_220 VDD VSS scs8hd_fill_2
XANTENNA__626__B x[27] VSS VDD scs8hd_diode_2
XFILLER_12_16 VSS VDD scs8hd_fill_1
XFILLER_12_27 VSS VDD scs8hd_decap_4
XFILLER_41_245 VSS VDD scs8hd_decap_8
X_340_ _336_/Y _337_/Y _693_/Q _337_/A _340_/X VSS VDD scs8hd_o22a_4
XANTENNA__552__A _552_/A VSS VDD scs8hd_diode_2
XFILLER_5_113 VDD VSS scs8hd_fill_2
XANTENNA__340__A2 _337_/Y VSS VDD scs8hd_diode_2
XANTENNA__695__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__628__B1 _624_/A VSS VDD scs8hd_diode_2
X_538_ _538_/A _538_/Y VSS VDD scs8hd_inv_8
X_607_ _602_/Y _603_/Y _683_/Q _603_/A _609_/B VSS VDD scs8hd_o22a_4
XANTENNA__646__RESETB _411_/X VSS VDD scs8hd_diode_2
X_469_ _469_/A _469_/X VSS VDD scs8hd_buf_1
XANTENNA__462__A _462_/A VSS VDD scs8hd_diode_2
XFILLER_23_245 VSS VDD scs8hd_decap_8
XFILLER_23_234 VDD VSS scs8hd_fill_2
XFILLER_23_223 VDD VSS scs8hd_fill_2
XFILLER_23_212 VDD VSS scs8hd_fill_2
XANTENNA__372__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_2_127 VSS VDD scs8hd_decap_4
XANTENNA__547__A _547_/A VSS VDD scs8hd_diode_2
XFILLER_9_39 VDD VSS scs8hd_fill_2
XFILLER_36_7 VDD VSS scs8hd_fill_2
XFILLER_1_160 VDD VSS scs8hd_fill_2
XFILLER_1_182 VSS VDD scs8hd_fill_1
XFILLER_20_215 VDD VSS scs8hd_fill_2
XFILLER_34_25 VDD VSS scs8hd_fill_2
XANTENNA__367__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_18_48 VSS VDD scs8hd_decap_12
XFILLER_34_69 VSS VDD scs8hd_decap_4
XFILLER_11_237 VSS VDD scs8hd_decap_6
XFILLER_24_91 VSS VDD scs8hd_fill_1
XFILLER_24_80 VSS VDD scs8hd_fill_1
XFILLER_6_241 VSS VDD scs8hd_decap_12
XFILLER_27_3 VSS VDD scs8hd_decap_4
XFILLER_37_123 VSS VDD scs8hd_decap_4
XFILLER_1_62 VDD VSS scs8hd_fill_2
XFILLER_1_73 VDD VSS scs8hd_fill_2
XANTENNA__470__A1 _466_/Y VSS VDD scs8hd_diode_2
XANTENNA__470__B2 _648_/Q VSS VDD scs8hd_diode_2
XFILLER_28_178 VDD VSS scs8hd_fill_2
XANTENNA__544__B _544_/B VSS VDD scs8hd_diode_2
XANTENNA__560__A _560_/A VSS VDD scs8hd_diode_2
XFILLER_10_93 VDD VSS scs8hd_fill_2
XFILLER_19_80 VDD VSS scs8hd_fill_2
XFILLER_19_91 VDD VSS scs8hd_fill_2
XFILLER_19_123 VDD VSS scs8hd_fill_2
XANTENNA__454__B x[3] VSS VDD scs8hd_diode_2
XANTENNA__443__B2 _442_/X VSS VDD scs8hd_diode_2
XFILLER_25_148 VSS VDD scs8hd_decap_3
XANTENNA__694__RESETB _353_/X VSS VDD scs8hd_diode_2
XFILLER_15_27 VDD VSS scs8hd_fill_2
XFILLER_33_192 VSS VDD scs8hd_fill_1
XFILLER_31_37 VDD VSS scs8hd_fill_2
XANTENNA__380__A _375_/A VSS VDD scs8hd_diode_2
X_640_ _648_/CLK _451_/X _640_/Q _418_/X VSS VDD scs8hd_dfrtp_4
X_571_ _567_/Y _568_/Y _673_/Q _676_/Q _573_/B VSS VDD scs8hd_o22a_4
XPHY_198 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__555__A _554_/X VSS VDD scs8hd_diode_2
XFILLER_24_181 VSS VDD scs8hd_decap_3
XPHY_187 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_110 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_121 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_132 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_143 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_154 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_16_159 VDD VSS scs8hd_fill_2
XPHY_165 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_176 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_1 VSS VDD scs8hd_decap_3
XANTENNA__465__A _462_/X VSS VDD scs8hd_diode_2
XFILLER_15_181 VDD VSS scs8hd_fill_2
XFILLER_26_37 VDD VSS scs8hd_fill_2
XANTENNA__375__A _375_/A VSS VDD scs8hd_diode_2
XFILLER_21_184 VSS VDD scs8hd_decap_3
X_485_ _481_/Y _482_/Y _649_/Q _652_/Q _485_/X VSS VDD scs8hd_o22a_4
X_554_ _547_/A x[17] _554_/X VSS VDD scs8hd_and2_4
X_623_ _623_/A _623_/B _688_/D VSS VDD scs8hd_xor2_4
XFILLER_12_151 VDD VSS scs8hd_fill_2
XANTENNA__642__RESETB _415_/X VSS VDD scs8hd_diode_2
XANTENNA__334__B1 _332_/X VSS VDD scs8hd_diode_2
XFILLER_5_158 VDD VSS scs8hd_fill_2
XANTENNA__628__B2 _625_/A VSS VDD scs8hd_diode_2
XANTENNA__628__A1 _624_/Y VSS VDD scs8hd_diode_2
X_537_ _534_/X _535_/X _537_/X VSS VDD scs8hd_xor2_4
XFILLER_32_224 VSS VDD scs8hd_decap_8
X_606_ _605_/X _609_/A VSS VDD scs8hd_buf_1
X_468_ _461_/A x[5] _469_/A VSS VDD scs8hd_and2_4
X_399_ _401_/A _399_/X VSS VDD scs8hd_buf_1
XANTENNA__564__B1 _671_/Q VSS VDD scs8hd_diode_2
XFILLER_4_84 VSS VDD scs8hd_decap_8
XANTENNA__547__B x[16] VSS VDD scs8hd_diode_2
XANTENNA__662__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_14_224 VSS VDD scs8hd_decap_3
XFILLER_13_82 VSS VDD scs8hd_decap_4
XANTENNA__563__A _563_/A VSS VDD scs8hd_diode_2
XFILLER_29_7 VSS VDD scs8hd_fill_1
XFILLER_38_90 VDD VSS scs8hd_fill_2
XANTENNA__473__A _473_/A VSS VDD scs8hd_diode_2
XFILLER_20_205 VSS VDD scs8hd_decap_4
XFILLER_18_16 VDD VSS scs8hd_fill_2
XFILLER_34_37 VSS VDD scs8hd_decap_8
XANTENNA__685__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__383__A _386_/A VSS VDD scs8hd_diode_2
XANTENNA__528__B1 _661_/Q VSS VDD scs8hd_diode_2
XFILLER_11_216 VDD VSS scs8hd_fill_2
XANTENNA__689__RESETB _360_/X VSS VDD scs8hd_diode_2
XANTENNA__558__A _558_/A VSS VDD scs8hd_diode_2
XFILLER_37_113 VSS VDD scs8hd_decap_4
XANTENNA__468__A _461_/A VSS VDD scs8hd_diode_2
XFILLER_1_85 VSS VDD scs8hd_decap_3
XANTENNA__470__A2 _467_/Y VSS VDD scs8hd_diode_2
XANTENNA__690__RESETB _357_/X VSS VDD scs8hd_diode_2
XFILLER_20_28 VSS VDD scs8hd_decap_3
XFILLER_29_48 VDD VSS scs8hd_fill_2
XFILLER_28_102 VDD VSS scs8hd_fill_2
XANTENNA__378__A _375_/A VSS VDD scs8hd_diode_2
XFILLER_3_245 VSS VDD scs8hd_decap_8
XFILLER_3_234 VDD VSS scs8hd_fill_2
XFILLER_10_83 VSS VDD scs8hd_decap_4
XFILLER_34_149 VSS VDD scs8hd_decap_4
XFILLER_34_127 VSS VDD scs8hd_decap_4
XFILLER_34_105 VSS VDD scs8hd_decap_8
XFILLER_19_168 VDD VSS scs8hd_fill_2
XFILLER_35_80 VDD VSS scs8hd_fill_2
XFILLER_40_119 VSS VDD scs8hd_decap_4
XFILLER_33_171 VDD VSS scs8hd_fill_2
XANTENNA__637__RESETB _421_/X VSS VDD scs8hd_diode_2
XFILLER_18_190 VDD VSS scs8hd_fill_2
XFILLER_31_27 VDD VSS scs8hd_fill_2
XFILLER_0_237 VSS VDD scs8hd_decap_8
XFILLER_0_226 VDD VSS scs8hd_fill_2
XPHY_100 VSS VDD scs8hd_tapvpwrvgnd_1
X_570_ _570_/A _570_/X VSS VDD scs8hd_buf_1
XPHY_199 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_188 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_177 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_111 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_122 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_133 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_144 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_155 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_166 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_2 VSS VDD scs8hd_decap_3
XANTENNA__465__B _465_/B VSS VDD scs8hd_diode_2
XFILLER_15_160 VDD VSS scs8hd_fill_2
XANTENNA__481__A _649_/Q VSS VDD scs8hd_diode_2
XFILLER_7_62 VDD VSS scs8hd_fill_2
XFILLER_7_95 VSS VDD scs8hd_fill_1
XFILLER_38_230 VSS VDD scs8hd_decap_6
XFILLER_42_48 VDD VSS scs8hd_fill_2
XFILLER_42_15 VSS VDD scs8hd_decap_12
XANTENNA__391__A _389_/A VSS VDD scs8hd_diode_2
XFILLER_13_108 VDD VSS scs8hd_fill_2
XFILLER_21_141 VSS VDD scs8hd_decap_3
XFILLER_21_174 VSS VDD scs8hd_fill_1
X_622_ _617_/Y _618_/Y _623_/A _623_/B _687_/D VSS VDD scs8hd_a2bb2o_4
X_484_ _483_/X _484_/X VSS VDD scs8hd_buf_1
X_553_ _553_/A _553_/Y VSS VDD scs8hd_inv_8
XANTENNA__566__A _566_/A VSS VDD scs8hd_diode_2
XFILLER_16_93 VDD VSS scs8hd_fill_2
XFILLER_8_101 VDD VSS scs8hd_fill_2
XFILLER_8_178 VDD VSS scs8hd_fill_2
XFILLER_12_163 VSS VDD scs8hd_decap_6
XANTENNA__476__A _476_/A VSS VDD scs8hd_diode_2
XFILLER_35_200 VDD VSS scs8hd_fill_2
XANTENNA__334__B2 _333_/X VSS VDD scs8hd_diode_2
XFILLER_41_236 VDD VSS scs8hd_fill_2
XFILLER_37_59 VDD VSS scs8hd_fill_2
XANTENNA__386__A _386_/A VSS VDD scs8hd_diode_2
XFILLER_5_137 VDD VSS scs8hd_fill_2
XANTENNA__628__A2 _625_/Y VSS VDD scs8hd_diode_2
X_605_ _605_/A x[24] _605_/X VSS VDD scs8hd_and2_4
X_536_ _531_/Y _532_/Y _534_/X _535_/X _536_/X VSS VDD scs8hd_a2bb2o_4
X_398_ _401_/A _398_/X VSS VDD scs8hd_buf_1
X_467_ _648_/Q _467_/Y VSS VDD scs8hd_inv_8
XANTENNA__564__B2 _560_/A VSS VDD scs8hd_diode_2
XANTENNA__564__A1 _559_/Y VSS VDD scs8hd_diode_2
XFILLER_4_74 VDD VSS scs8hd_fill_2
XFILLER_4_41 VSS VDD scs8hd_decap_4
XFILLER_4_30 VSS VDD scs8hd_fill_1
XANTENNA__457__A2N _453_/Y VSS VDD scs8hd_diode_2
XANTENNA__685__RESETB _364_/X VSS VDD scs8hd_diode_2
XFILLER_1_184 VSS VDD scs8hd_decap_4
X_519_ _547_/A x[12] _519_/X VSS VDD scs8hd_and2_4
XFILLER_20_239 VSS VDD scs8hd_decap_12
XANTENNA__528__A1 _524_/Y VSS VDD scs8hd_diode_2
XANTENNA__528__B2 _664_/Q VSS VDD scs8hd_diode_2
XANTENNA__464__B1 _462_/X VSS VDD scs8hd_diode_2
XANTENNA__558__B _558_/B VSS VDD scs8hd_diode_2
XFILLER_24_93 VSS VDD scs8hd_decap_6
XANTENNA__574__A _574_/A VSS VDD scs8hd_diode_2
XFILLER_10_250 VSS VDD scs8hd_decap_3
XFILLER_6_221 VDD VSS scs8hd_fill_2
XANTENNA__468__B x[5] VSS VDD scs8hd_diode_2
XFILLER_1_53 VSS VDD scs8hd_decap_4
XANTENNA__622__A2N _618_/Y VSS VDD scs8hd_diode_2
XANTENNA__484__A _483_/X VSS VDD scs8hd_diode_2
XANTENNA__634__D _634_/D VSS VDD scs8hd_diode_2
XANTENNA__652__CLK _651_/CLK VSS VDD scs8hd_diode_2
XANTENNA__633__RESETB _425_/X VSS VDD scs8hd_diode_2
XFILLER_36_180 VDD VSS scs8hd_fill_2
XFILLER_28_147 VDD VSS scs8hd_fill_2
XANTENNA__394__A _389_/A VSS VDD scs8hd_diode_2
XANTENNA__569__A _597_/A VSS VDD scs8hd_diode_2
XFILLER_19_103 VSS VDD scs8hd_decap_4
XFILLER_19_114 VSS VDD scs8hd_decap_4
XFILLER_42_161 VSS VDD scs8hd_decap_8
XANTENNA__675__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_32_3 VDD VSS scs8hd_fill_2
XFILLER_25_128 VDD VSS scs8hd_fill_2
XFILLER_25_117 VSS VDD scs8hd_decap_4
XANTENNA__600__B1 _598_/X VSS VDD scs8hd_diode_2
XANTENNA__389__A _389_/A VSS VDD scs8hd_diode_2
XFILLER_0_249 VSS VDD scs8hd_decap_4
XPHY_101 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_112 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_123 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_134 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_16_139 VSS VDD scs8hd_decap_6
XPHY_189 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_178 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_145 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_156 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_167 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_11_8 VDD VSS scs8hd_fill_2
XFILLER_30_131 VDD VSS scs8hd_fill_2
XPHY_3 VSS VDD scs8hd_decap_3
XFILLER_30_186 VDD VSS scs8hd_fill_2
XFILLER_30_175 VDD VSS scs8hd_fill_2
XFILLER_7_52 VSS VDD scs8hd_decap_4
XFILLER_26_17 VDD VSS scs8hd_fill_2
XFILLER_42_27 VSS VDD scs8hd_decap_4
XFILLER_21_120 VDD VSS scs8hd_fill_2
X_621_ _617_/Y _618_/Y _687_/Q _690_/Q _623_/B VSS VDD scs8hd_o22a_4
XANTENNA__582__A _582_/A VSS VDD scs8hd_diode_2
X_483_ _476_/A x[7] _483_/X VSS VDD scs8hd_and2_4
X_552_ _552_/A _552_/Y VSS VDD scs8hd_inv_8
XANTENNA__566__B _566_/B VSS VDD scs8hd_diode_2
XFILLER_16_61 VDD VSS scs8hd_fill_2
XFILLER_32_93 VDD VSS scs8hd_fill_2
XFILLER_8_113 VSS VDD scs8hd_fill_1
XFILLER_12_175 VSS VDD scs8hd_fill_1
XANTENNA__476__B x[6] VSS VDD scs8hd_diode_2
XFILLER_35_245 VSS VDD scs8hd_decap_8
XANTENNA__642__D _458_/X VSS VDD scs8hd_diode_2
XFILLER_12_19 VDD VSS scs8hd_fill_2
XFILLER_37_38 VSS VDD scs8hd_fill_1
XFILLER_26_212 VDD VSS scs8hd_fill_2
XFILLER_5_127 VSS VDD scs8hd_decap_3
XANTENNA__681__RESETB _369_/X VSS VDD scs8hd_diode_2
X_535_ _531_/Y _532_/Y _663_/Q _666_/Q _535_/X VSS VDD scs8hd_o22a_4
XFILLER_27_82 VSS VDD scs8hd_decap_3
X_604_ y _605_/A VSS VDD scs8hd_buf_1
XANTENNA__577__A _577_/A VSS VDD scs8hd_diode_2
XFILLER_17_245 VDD VSS scs8hd_fill_2
XFILLER_32_215 VDD VSS scs8hd_fill_2
X_466_ _645_/Q _466_/Y VSS VDD scs8hd_inv_8
XANTENNA__564__A2 _560_/Y VSS VDD scs8hd_diode_2
X_397_ _401_/A _397_/X VSS VDD scs8hd_buf_1
XFILLER_4_193 VDD VSS scs8hd_fill_2
XANTENNA__487__A _484_/X VSS VDD scs8hd_diode_2
XANTENNA__637__D _443_/X VSS VDD scs8hd_diode_2
XANTENNA__397__A _401_/A VSS VDD scs8hd_diode_2
XANTENNA__457__A1N _452_/Y VSS VDD scs8hd_diode_2
XFILLER_13_40 VSS VDD scs8hd_decap_4
XFILLER_13_51 VDD VSS scs8hd_fill_2
XFILLER_14_215 VDD VSS scs8hd_fill_2
XFILLER_13_62 VDD VSS scs8hd_fill_2
XFILLER_1_174 VDD VSS scs8hd_fill_2
X_518_ _518_/A _547_/A VSS VDD scs8hd_buf_1
X_449_ _445_/Y _446_/Y _445_/A _446_/A _449_/X VSS VDD scs8hd_o22a_4
XFILLER_9_241 VSS VDD scs8hd_decap_3
XFILLER_18_29 VDD VSS scs8hd_fill_2
XANTENNA__528__A2 _525_/Y VSS VDD scs8hd_diode_2
XFILLER_11_229 VDD VSS scs8hd_fill_2
XANTENNA__464__B2 _465_/B VSS VDD scs8hd_diode_2
XANTENNA__590__A _597_/A VSS VDD scs8hd_diode_2
XFILLER_24_83 VSS VDD scs8hd_decap_8
XFILLER_24_72 VSS VDD scs8hd_decap_8
XFILLER_24_61 VSS VDD scs8hd_decap_4
XFILLER_40_93 VSS VDD scs8hd_decap_4
XANTENNA__622__A1N _617_/Y VSS VDD scs8hd_diode_2
XFILLER_1_43 VSS VDD scs8hd_fill_1
XANTENNA__650__D _487_/X VSS VDD scs8hd_diode_2
XFILLER_29_39 VSS VDD scs8hd_decap_3
XFILLER_28_137 VSS VDD scs8hd_fill_1
XFILLER_3_214 VDD VSS scs8hd_fill_2
XFILLER_10_30 VSS VDD scs8hd_fill_1
XANTENNA__437__A1 _635_/Q VSS VDD scs8hd_diode_2
XANTENNA__569__B x[19] VSS VDD scs8hd_diode_2
XFILLER_19_137 VSS VDD scs8hd_fill_1
XFILLER_34_118 VDD VSS scs8hd_fill_2
XFILLER_27_181 VDD VSS scs8hd_fill_2
XFILLER_25_3 VDD VSS scs8hd_fill_2
XANTENNA__495__A _653_/Q VSS VDD scs8hd_diode_2
XANTENNA__600__B2 _601_/B VSS VDD scs8hd_diode_2
XFILLER_33_195 VDD VSS scs8hd_fill_2
XFILLER_33_184 VDD VSS scs8hd_fill_2
XANTENNA__645__D _471_/X VSS VDD scs8hd_diode_2
XFILLER_24_173 VSS VDD scs8hd_decap_8
XPHY_102 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_113 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_124 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_135 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_146 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_157 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_179 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_168 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_21_40 VDD VSS scs8hd_fill_2
XFILLER_21_51 VDD VSS scs8hd_fill_2
XFILLER_21_62 VDD VSS scs8hd_fill_2
XFILLER_30_165 VSS VDD scs8hd_decap_3
XFILLER_30_154 VDD VSS scs8hd_fill_2
XFILLER_30_143 VDD VSS scs8hd_fill_2
XPHY_4 VSS VDD scs8hd_decap_3
XANTENNA__642__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_15_140 VSS VDD scs8hd_fill_1
XFILLER_15_184 VDD VSS scs8hd_fill_2
XANTENNA__676__RESETB _376_/X VSS VDD scs8hd_diode_2
XFILLER_30_198 VDD VSS scs8hd_fill_2
XFILLER_7_42 VSS VDD scs8hd_decap_3
XANTENNA__585__B1 _581_/A VSS VDD scs8hd_diode_2
XFILLER_26_29 VDD VSS scs8hd_fill_2
XFILLER_21_110 VDD VSS scs8hd_fill_2
XFILLER_21_154 VDD VSS scs8hd_fill_2
X_551_ _548_/X _551_/B _551_/X VSS VDD scs8hd_xor2_4
XANTENNA__665__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_29_243 VSS VDD scs8hd_fill_1
X_620_ _620_/A _623_/A VSS VDD scs8hd_buf_1
X_482_ _652_/Q _482_/Y VSS VDD scs8hd_inv_8
XFILLER_12_154 VDD VSS scs8hd_fill_2
XFILLER_12_187 VDD VSS scs8hd_fill_2
XFILLER_8_147 VDD VSS scs8hd_fill_2
XFILLER_12_198 VDD VSS scs8hd_fill_2
XANTENNA__500__B1 _498_/X VSS VDD scs8hd_diode_2
XFILLER_35_213 VSS VDD scs8hd_decap_4
XANTENNA__688__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_41_227 VDD VSS scs8hd_fill_2
XFILLER_41_216 VDD VSS scs8hd_fill_2
XFILLER_5_117 VSS VDD scs8hd_decap_4
XANTENNA__549__B1 _545_/A VSS VDD scs8hd_diode_2
X_534_ _533_/X _534_/X VSS VDD scs8hd_buf_1
X_603_ _603_/A _603_/Y VSS VDD scs8hd_inv_8
X_465_ _462_/X _465_/B _465_/X VSS VDD scs8hd_xor2_4
XFILLER_17_213 VSS VDD scs8hd_decap_3
X_396_ _401_/A _396_/X VSS VDD scs8hd_buf_1
XFILLER_4_32 VDD VSS scs8hd_fill_2
XANTENNA__487__B _485_/X VSS VDD scs8hd_diode_2
XFILLER_4_98 VSS VDD scs8hd_decap_12
XANTENNA__653__D _653_/D VSS VDD scs8hd_diode_2
XFILLER_23_238 VDD VSS scs8hd_fill_2
XFILLER_23_227 VSS VDD scs8hd_decap_4
XFILLER_1_120 VDD VSS scs8hd_fill_2
XFILLER_38_93 VDD VSS scs8hd_fill_2
XANTENNA__588__A _679_/Q VSS VDD scs8hd_diode_2
XFILLER_1_164 VSS VDD scs8hd_decap_4
X_517_ _662_/Q _517_/Y VSS VDD scs8hd_inv_8
X_448_ _448_/A _451_/A VSS VDD scs8hd_buf_1
X_379_ _375_/A _379_/X VSS VDD scs8hd_buf_1
XANTENNA__498__A _497_/X VSS VDD scs8hd_diode_2
XANTENNA__648__D _480_/X VSS VDD scs8hd_diode_2
XFILLER_34_29 VDD VSS scs8hd_fill_2
XFILLER_1_8 VDD VSS scs8hd_fill_2
XFILLER_39_190 VDD VSS scs8hd_fill_2
XANTENNA__590__B x[22] VSS VDD scs8hd_diode_2
XFILLER_6_212 VDD VSS scs8hd_fill_2
XFILLER_37_127 VSS VDD scs8hd_fill_1
XFILLER_1_77 VSS VDD scs8hd_decap_8
XFILLER_1_99 VDD VSS scs8hd_fill_2
XFILLER_28_116 VSS VDD scs8hd_decap_8
XFILLER_36_171 VSS VDD scs8hd_decap_6
XFILLER_10_53 VDD VSS scs8hd_fill_2
XFILLER_10_64 VDD VSS scs8hd_fill_2
XFILLER_10_75 VDD VSS scs8hd_fill_2
XANTENNA__437__A2 _435_/X VSS VDD scs8hd_diode_2
XFILLER_27_171 VSS VDD scs8hd_decap_4
XFILLER_19_62 VSS VDD scs8hd_decap_4
XFILLER_19_84 VSS VDD scs8hd_decap_4
XFILLER_19_95 VDD VSS scs8hd_fill_2
XANTENNA__672__RESETB _380_/X VSS VDD scs8hd_diode_2
XFILLER_18_3 VDD VSS scs8hd_fill_2
XFILLER_33_163 VDD VSS scs8hd_fill_2
XFILLER_18_182 VDD VSS scs8hd_fill_2
XANTENNA__661__D _661_/D VSS VDD scs8hd_diode_2
XFILLER_0_218 VDD VSS scs8hd_fill_2
XPHY_103 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_114 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_125 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_136 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_147 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_158 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_169 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__596__A _684_/Q VSS VDD scs8hd_diode_2
X_696_ _681_/CLK _349_/X _337_/A _350_/X VSS VDD scs8hd_dfrtp_4
XPHY_5 VSS VDD scs8hd_decap_3
XFILLER_15_152 VDD VSS scs8hd_fill_2
XFILLER_7_87 VDD VSS scs8hd_fill_2
XFILLER_38_222 VDD VSS scs8hd_fill_2
XANTENNA__585__B2 _582_/A VSS VDD scs8hd_diode_2
XANTENNA__585__A1 _581_/Y VSS VDD scs8hd_diode_2
XANTENNA__656__D _508_/X VSS VDD scs8hd_diode_2
XFILLER_21_177 VDD VSS scs8hd_fill_2
X_550_ _545_/Y _546_/Y _548_/X _551_/B _550_/X VSS VDD scs8hd_a2bb2o_4
X_481_ _649_/Q _481_/Y VSS VDD scs8hd_inv_8
XFILLER_29_233 VDD VSS scs8hd_fill_2
XFILLER_29_222 VDD VSS scs8hd_fill_2
XFILLER_8_137 VSS VDD scs8hd_decap_4
XANTENNA__500__B2 _501_/B VSS VDD scs8hd_diode_2
XFILLER_35_236 VDD VSS scs8hd_fill_2
X_679_ _667_/CLK _593_/X _679_/Q _371_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_181 VDD VSS scs8hd_fill_2
X_602_ _683_/Q _602_/Y VSS VDD scs8hd_inv_8
X_533_ _547_/A x[14] _533_/X VSS VDD scs8hd_and2_4
XANTENNA__549__A1 _545_/Y VSS VDD scs8hd_diode_2
XANTENNA__549__B2 _546_/A VSS VDD scs8hd_diode_2
XFILLER_32_206 VSS VDD scs8hd_decap_8
XFILLER_27_73 VSS VDD scs8hd_decap_6
XFILLER_27_62 VDD VSS scs8hd_fill_2
XFILLER_27_51 VDD VSS scs8hd_fill_2
X_464_ _459_/Y _460_/Y _462_/X _465_/B _643_/D VSS VDD scs8hd_a2bb2o_4
XFILLER_17_236 VDD VSS scs8hd_fill_2
X_395_ _402_/A _401_/A VSS VDD scs8hd_buf_1
XANTENNA__485__B1 _649_/Q VSS VDD scs8hd_diode_2
XFILLER_4_184 VDD VSS scs8hd_fill_2
XFILLER_4_151 VDD VSS scs8hd_fill_2
XFILLER_4_66 VDD VSS scs8hd_fill_2
XFILLER_4_22 VDD VSS scs8hd_fill_2
XFILLER_4_11 VDD VSS scs8hd_fill_2
XANTENNA__655__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_14_206 VSS VDD scs8hd_decap_8
XFILLER_13_86 VSS VDD scs8hd_fill_1
XFILLER_1_132 VDD VSS scs8hd_fill_2
X_516_ _516_/A _516_/Y VSS VDD scs8hd_inv_8
X_447_ _461_/A x[2] _448_/A VSS VDD scs8hd_and2_4
X_378_ _375_/A _378_/X VSS VDD scs8hd_buf_1
XFILLER_20_209 VSS VDD scs8hd_fill_1
XANTENNA__678__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__667__RESETB _386_/X VSS VDD scs8hd_diode_2
XANTENNA__664__D _537_/X VSS VDD scs8hd_diode_2
XFILLER_11_209 VSS VDD scs8hd_decap_4
XANTENNA__449__B1 _445_/A VSS VDD scs8hd_diode_2
XFILLER_39_180 VSS VDD scs8hd_decap_3
XANTENNA__621__B1 _687_/Q VSS VDD scs8hd_diode_2
XFILLER_40_84 VDD VSS scs8hd_fill_2
XFILLER_40_73 VSS VDD scs8hd_decap_4
XFILLER_6_202 VSS VDD scs8hd_fill_1
XFILLER_10_220 VDD VSS scs8hd_fill_2
XFILLER_10_231 VDD VSS scs8hd_fill_2
XFILLER_10_242 VSS VDD scs8hd_decap_8
XFILLER_1_23 VDD VSS scs8hd_fill_2
XFILLER_37_117 VSS VDD scs8hd_fill_1
XFILLER_1_34 VSS VDD scs8hd_decap_3
XFILLER_28_106 VDD VSS scs8hd_fill_2
XANTENNA__659__D _522_/X VSS VDD scs8hd_diode_2
XANTENNA__493__A2N _489_/Y VSS VDD scs8hd_diode_2
XFILLER_3_238 VSS VDD scs8hd_decap_6
XFILLER_10_32 VDD VSS scs8hd_fill_2
XFILLER_10_87 VSS VDD scs8hd_fill_1
XFILLER_19_41 VSS VDD scs8hd_decap_4
XFILLER_42_142 VDD VSS scs8hd_fill_2
XFILLER_35_84 VDD VSS scs8hd_fill_2
XFILLER_35_62 VSS VDD scs8hd_decap_12
XFILLER_33_175 VSS VDD scs8hd_decap_8
XFILLER_25_109 VDD VSS scs8hd_fill_2
XFILLER_24_197 VDD VSS scs8hd_fill_2
XFILLER_24_186 VDD VSS scs8hd_fill_2
XPHY_104 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_115 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_126 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_137 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_148 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_159 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_6 VSS VDD scs8hd_decap_3
X_695_ _681_/CLK _348_/X _343_/A _357_/A VSS VDD scs8hd_dfrtp_4
XFILLER_15_164 VDD VSS scs8hd_fill_2
XFILLER_15_175 VSS VDD scs8hd_decap_4
XFILLER_30_3 VDD VSS scs8hd_fill_2
XFILLER_7_99 VDD VSS scs8hd_fill_2
XFILLER_38_245 VSS VDD scs8hd_decap_8
XANTENNA__585__A2 _582_/Y VSS VDD scs8hd_diode_2
XANTENNA__672__D _672_/D VSS VDD scs8hd_diode_2
XFILLER_21_123 VDD VSS scs8hd_fill_2
XFILLER_21_189 VDD VSS scs8hd_fill_2
XFILLER_29_245 VSS VDD scs8hd_decap_8
X_480_ _477_/X _480_/B _480_/X VSS VDD scs8hd_xor2_4
XFILLER_16_20 VDD VSS scs8hd_fill_2
XFILLER_32_85 VSS VDD scs8hd_decap_3
XFILLER_32_52 VDD VSS scs8hd_fill_2
XFILLER_8_105 VSS VDD scs8hd_decap_8
XFILLER_12_178 VDD VSS scs8hd_fill_2
XFILLER_35_204 VDD VSS scs8hd_fill_2
XANTENNA__400__A _401_/A VSS VDD scs8hd_diode_2
X_678_ _667_/CLK _587_/X _678_/Q _372_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_171 VSS VDD scs8hd_decap_4
XANTENNA__667__D _550_/X VSS VDD scs8hd_diode_2
XFILLER_26_237 VSS VDD scs8hd_decap_12
XFILLER_26_215 VDD VSS scs8hd_fill_2
X_601_ _598_/X _601_/B _601_/X VSS VDD scs8hd_xor2_4
XFILLER_40_240 VSS VDD scs8hd_decap_12
XANTENNA__549__A2 _546_/Y VSS VDD scs8hd_diode_2
X_532_ _666_/Q _532_/Y VSS VDD scs8hd_inv_8
X_394_ _389_/A _394_/X VSS VDD scs8hd_buf_1
X_463_ _459_/Y _460_/Y _643_/Q _460_/A _465_/B VSS VDD scs8hd_o22a_4
X_CTS_root clk _CTS_root/X VSS VDD scs8hd_clkbuf_16
XANTENNA__485__B2 _652_/Q VSS VDD scs8hd_diode_2
XANTENNA__485__A1 _481_/Y VSS VDD scs8hd_diode_2
XFILLER_4_78 VSS VDD scs8hd_decap_3
XFILLER_4_45 VSS VDD scs8hd_fill_1
XANTENNA__663__RESETB _391_/X VSS VDD scs8hd_diode_2
XFILLER_22_251 VDD VSS scs8hd_fill_2
XFILLER_14_229 VSS VDD scs8hd_decap_4
XFILLER_1_188 VSS VDD scs8hd_fill_1
XFILLER_8_3 VDD VSS scs8hd_fill_2
XFILLER_38_84 VSS VDD scs8hd_decap_4
XFILLER_38_73 VSS VDD scs8hd_decap_8
XFILLER_38_62 VDD VSS scs8hd_fill_2
X_515_ _515_/A _513_/X _515_/X VSS VDD scs8hd_xor2_4
X_377_ _375_/A _377_/X VSS VDD scs8hd_buf_1
XFILLER_9_211 VDD VSS scs8hd_fill_2
X_446_ _446_/A _446_/Y VSS VDD scs8hd_inv_8
XFILLER_13_240 VSS VDD scs8hd_decap_4
XANTENNA__680__D _680_/D VSS VDD scs8hd_diode_2
XANTENNA__449__B2 _446_/A VSS VDD scs8hd_diode_2
XANTENNA__449__A1 _445_/Y VSS VDD scs8hd_diode_2
XANTENNA__621__B2 _690_/Q VSS VDD scs8hd_diode_2
XANTENNA__621__A1 _617_/Y VSS VDD scs8hd_diode_2
XFILLER_10_210 VSS VDD scs8hd_decap_4
XANTENNA__615__A2N _611_/Y VSS VDD scs8hd_diode_2
XFILLER_40_52 VSS VDD scs8hd_decap_4
XFILLER_27_9 VDD VSS scs8hd_fill_2
XANTENNA__645__CLK _648_/CLK VSS VDD scs8hd_diode_2
X_429_ _518_/A _461_/A VSS VDD scs8hd_buf_1
XANTENNA__493__A1N _488_/Y VSS VDD scs8hd_diode_2
XANTENNA__675__D _579_/X VSS VDD scs8hd_diode_2
XFILLER_10_11 VDD VSS scs8hd_fill_2
XFILLER_10_22 VDD VSS scs8hd_fill_2
XFILLER_19_20 VDD VSS scs8hd_fill_2
XFILLER_19_53 VSS VDD scs8hd_decap_4
XFILLER_19_107 VSS VDD scs8hd_fill_1
XFILLER_42_154 VSS VDD scs8hd_fill_1
XANTENNA__668__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_35_74 VSS VDD scs8hd_decap_4
XFILLER_27_184 VDD VSS scs8hd_fill_2
XFILLER_42_187 VSS VDD scs8hd_decap_12
XFILLER_32_7 VSS VDD scs8hd_decap_3
XANTENNA__403__A _405_/A VSS VDD scs8hd_diode_2
XFILLER_18_151 VDD VSS scs8hd_fill_2
XFILLER_18_195 VDD VSS scs8hd_fill_2
XANTENNA__521__B1 _516_/A VSS VDD scs8hd_diode_2
XFILLER_0_209 VDD VSS scs8hd_fill_2
XPHY_105 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_116 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_24_154 VSS VDD scs8hd_decap_6
XPHY_127 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_138 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_149 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_21_87 VDD VSS scs8hd_fill_2
X_694_ _681_/CLK _694_/D _694_/Q _353_/X VSS VDD scs8hd_dfrtp_4
XFILLER_30_135 VSS VDD scs8hd_decap_8
XFILLER_30_102 VDD VSS scs8hd_fill_2
XPHY_7 VSS VDD scs8hd_decap_3
XFILLER_15_132 VDD VSS scs8hd_fill_2
XFILLER_15_143 VDD VSS scs8hd_fill_2
XANTENNA__579__B1 _580_/A VSS VDD scs8hd_diode_2
XFILLER_30_179 VSS VDD scs8hd_decap_4
XFILLER_7_12 VDD VSS scs8hd_fill_2
XFILLER_7_56 VSS VDD scs8hd_fill_1
XFILLER_7_78 VDD VSS scs8hd_fill_2
XFILLER_38_202 VDD VSS scs8hd_fill_2
XFILLER_23_3 VSS VDD scs8hd_decap_4
XFILLER_21_102 VDD VSS scs8hd_fill_2
XFILLER_21_146 VDD VSS scs8hd_fill_2
XFILLER_12_113 VSS VDD scs8hd_decap_8
XFILLER_16_32 VDD VSS scs8hd_fill_2
XFILLER_16_65 VSS VDD scs8hd_decap_4
XFILLER_16_98 VSS VDD scs8hd_decap_3
XANTENNA__658__RESETB _397_/X VSS VDD scs8hd_diode_2
X_677_ _667_/CLK _586_/X _581_/A _375_/X VSS VDD scs8hd_dfrtp_4
XFILLER_41_208 VSS VDD scs8hd_decap_6
XFILLER_26_249 VSS VDD scs8hd_decap_4
XANTENNA__683__D _683_/D VSS VDD scs8hd_diode_2
XFILLER_5_109 VDD VSS scs8hd_fill_2
XANTENNA__501__A _498_/X VSS VDD scs8hd_diode_2
X_600_ _595_/Y _596_/Y _598_/X _601_/B _600_/X VSS VDD scs8hd_a2bb2o_4
X_531_ _663_/Q _531_/Y VSS VDD scs8hd_inv_8
XFILLER_17_249 VSS VDD scs8hd_decap_4
XFILLER_40_252 VSS VDD scs8hd_fill_1
X_393_ _389_/A _393_/X VSS VDD scs8hd_buf_1
X_462_ _462_/A _462_/X VSS VDD scs8hd_buf_1
XFILLER_4_120 VSS VDD scs8hd_fill_1
XANTENNA__485__A2 _482_/Y VSS VDD scs8hd_diode_2
XFILLER_4_197 VSS VDD scs8hd_decap_8
XANTENNA__411__A _410_/A VSS VDD scs8hd_diode_2
XFILLER_23_208 VDD VSS scs8hd_fill_2
XANTENNA__678__D _587_/X VSS VDD scs8hd_diode_2
XFILLER_13_11 VDD VSS scs8hd_fill_2
XFILLER_13_44 VSS VDD scs8hd_fill_1
XFILLER_13_55 VDD VSS scs8hd_fill_2
XFILLER_1_178 VSS VDD scs8hd_decap_4
XFILLER_1_123 VDD VSS scs8hd_fill_2
X_514_ _509_/Y _510_/Y _515_/A _513_/X _514_/X VSS VDD scs8hd_a2bb2o_4
XANTENNA__406__A _405_/A VSS VDD scs8hd_diode_2
X_445_ _445_/A _445_/Y VSS VDD scs8hd_inv_8
XFILLER_9_245 VSS VDD scs8hd_decap_8
X_376_ _375_/A _376_/X VSS VDD scs8hd_buf_1
XANTENNA__449__A2 _446_/Y VSS VDD scs8hd_diode_2
XANTENNA__621__A2 _618_/Y VSS VDD scs8hd_diode_2
XANTENNA__615__A1N _610_/Y VSS VDD scs8hd_diode_2
XFILLER_24_65 VSS VDD scs8hd_fill_1
XFILLER_24_32 VDD VSS scs8hd_fill_2
XFILLER_24_21 VDD VSS scs8hd_fill_2
XFILLER_6_215 VSS VDD scs8hd_decap_4
XFILLER_6_237 VDD VSS scs8hd_fill_2
X_428_ y _518_/A VSS VDD scs8hd_buf_1
X_359_ _366_/A _363_/A VSS VDD scs8hd_buf_1
XFILLER_36_163 VSS VDD scs8hd_decap_4
XFILLER_36_130 VDD VSS scs8hd_fill_2
XANTENNA__691__D _691_/D VSS VDD scs8hd_diode_2
XFILLER_10_45 VSS VDD scs8hd_decap_6
XFILLER_19_76 VDD VSS scs8hd_fill_2
XFILLER_42_122 VDD VSS scs8hd_fill_2
XFILLER_35_42 VDD VSS scs8hd_fill_2
XFILLER_27_130 VDD VSS scs8hd_fill_2
XFILLER_42_199 VSS VDD scs8hd_decap_12
XFILLER_2_240 VSS VDD scs8hd_decap_12
XFILLER_33_111 VSS VDD scs8hd_decap_8
XFILLER_33_100 VSS VDD scs8hd_decap_4
XFILLER_18_163 VDD VSS scs8hd_fill_2
XFILLER_33_199 VDD VSS scs8hd_fill_2
XFILLER_33_188 VSS VDD scs8hd_decap_4
XFILLER_33_133 VSS VDD scs8hd_decap_3
XANTENNA__521__A1 _516_/Y VSS VDD scs8hd_diode_2
XANTENNA__521__B2 _662_/Q VSS VDD scs8hd_diode_2
XANTENNA__686__D _686_/D VSS VDD scs8hd_diode_2
XFILLER_24_111 VSS VDD scs8hd_decap_12
XPHY_106 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_117 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_128 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_139 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__504__A _476_/A VSS VDD scs8hd_diode_2
XFILLER_21_44 VSS VDD scs8hd_decap_4
XFILLER_21_55 VDD VSS scs8hd_fill_2
XANTENNA__654__RESETB _401_/X VSS VDD scs8hd_diode_2
XANTENNA__635__CLK _648_/CLK VSS VDD scs8hd_diode_2
X_693_ _681_/CLK _341_/X _693_/Q _354_/X VSS VDD scs8hd_dfrtp_4
XFILLER_15_100 VSS VDD scs8hd_decap_4
XANTENNA__579__B2 _578_/X VSS VDD scs8hd_diode_2
XFILLER_30_147 VSS VDD scs8hd_decap_6
XPHY_8 VSS VDD scs8hd_decap_3
XANTENNA__414__A _410_/A VSS VDD scs8hd_diode_2
XFILLER_16_3 VDD VSS scs8hd_fill_2
XANTENNA__658__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_21_114 VSS VDD scs8hd_decap_4
XFILLER_12_136 VSS VDD scs8hd_decap_12
XFILLER_32_32 VSS VDD scs8hd_decap_4
XFILLER_20_191 VSS VDD scs8hd_decap_4
XFILLER_35_217 VSS VDD scs8hd_fill_1
XANTENNA__409__A _402_/A VSS VDD scs8hd_diode_2
X_676_ _667_/CLK _580_/X _676_/Q _376_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__450__A2N _446_/Y VSS VDD scs8hd_diode_2
XFILLER_7_184 VSS VDD scs8hd_decap_4
XANTENNA__479__B1 _477_/X VSS VDD scs8hd_diode_2
XANTENNA__501__B _501_/B VSS VDD scs8hd_diode_2
X_530_ _527_/X _528_/X _662_/D VSS VDD scs8hd_xor2_4
XFILLER_27_87 VDD VSS scs8hd_fill_2
X_461_ _461_/A x[4] _462_/A VSS VDD scs8hd_and2_4
X_392_ _389_/A _392_/X VSS VDD scs8hd_buf_1
XFILLER_4_154 VDD VSS scs8hd_fill_2
XFILLER_4_132 VDD VSS scs8hd_fill_2
XFILLER_4_110 VSS VDD scs8hd_fill_1
X_659_ _651_/CLK _522_/X _516_/A _396_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__602__A _683_/Q VSS VDD scs8hd_diode_2
XANTENNA__694__D _694_/D VSS VDD scs8hd_diode_2
XFILLER_1_113 VSS VDD scs8hd_decap_4
XFILLER_13_78 VDD VSS scs8hd_fill_2
XFILLER_13_89 VDD VSS scs8hd_fill_2
XANTENNA__512__A _512_/A VSS VDD scs8hd_diode_2
X_513_ _509_/Y _510_/Y _657_/Q _660_/Q _513_/X VSS VDD scs8hd_o22a_4
X_444_ _441_/X _442_/X _444_/X VSS VDD scs8hd_xor2_4
X_375_ _375_/A _375_/X VSS VDD scs8hd_buf_1
XFILLER_9_202 VSS VDD scs8hd_decap_3
XFILLER_9_235 VSS VDD scs8hd_decap_4
XANTENNA__422__A _417_/A VSS VDD scs8hd_diode_2
XANTENNA__615__B1 _616_/A VSS VDD scs8hd_diode_2
XANTENNA__332__A _331_/X VSS VDD scs8hd_diode_2
XANTENNA__689__D _629_/X VSS VDD scs8hd_diode_2
XFILLER_39_194 VDD VSS scs8hd_fill_2
XFILLER_39_172 VDD VSS scs8hd_fill_2
XFILLER_40_32 VSS VDD scs8hd_decap_4
XFILLER_6_205 VSS VDD scs8hd_decap_4
XFILLER_1_59 VDD VSS scs8hd_fill_2
XANTENNA__649__RESETB _407_/X VSS VDD scs8hd_diode_2
X_427_ _638_/Q _427_/Y VSS VDD scs8hd_inv_8
X_358_ _373_/A _366_/A VSS VDD scs8hd_buf_1
XANTENNA__417__A _417_/A VSS VDD scs8hd_diode_2
XANTENNA__691__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_3_208 VSS VDD scs8hd_decap_4
XFILLER_10_68 VSS VDD scs8hd_decap_4
XFILLER_10_79 VDD VSS scs8hd_fill_2
XFILLER_27_120 VDD VSS scs8hd_fill_2
XFILLER_19_66 VSS VDD scs8hd_fill_1
XFILLER_19_88 VSS VDD scs8hd_fill_1
XFILLER_19_99 VDD VSS scs8hd_fill_2
XFILLER_42_178 VSS VDD scs8hd_decap_8
XFILLER_42_156 VDD VSS scs8hd_fill_2
XANTENNA__650__RESETB _406_/X VSS VDD scs8hd_diode_2
XFILLER_2_252 VSS VDD scs8hd_fill_1
XFILLER_33_123 VDD VSS scs8hd_fill_2
XANTENNA__557__A2N _553_/Y VSS VDD scs8hd_diode_2
XFILLER_18_142 VDD VSS scs8hd_fill_2
XFILLER_18_186 VDD VSS scs8hd_fill_2
XFILLER_33_167 VDD VSS scs8hd_fill_2
XANTENNA__521__A2 _517_/Y VSS VDD scs8hd_diode_2
XFILLER_2_91 VSS VDD scs8hd_fill_1
XANTENNA__610__A _685_/Q VSS VDD scs8hd_diode_2
XPHY_107 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_118 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_129 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__504__B x[10] VSS VDD scs8hd_diode_2
XFILLER_21_12 VSS VDD scs8hd_fill_1
XANTENNA__520__A _519_/X VSS VDD scs8hd_diode_2
XPHY_9 VSS VDD scs8hd_decap_3
X_692_ _681_/CLK _692_/D _625_/A _355_/X VSS VDD scs8hd_dfrtp_4
XFILLER_15_123 VDD VSS scs8hd_fill_2
XFILLER_15_156 VDD VSS scs8hd_fill_2
XFILLER_38_226 VDD VSS scs8hd_fill_2
XFILLER_38_215 VSS VDD scs8hd_decap_4
XANTENNA__430__A _461_/A VSS VDD scs8hd_diode_2
XANTENNA__605__A _605_/A VSS VDD scs8hd_diode_2
XFILLER_29_237 VSS VDD scs8hd_decap_6
XFILLER_29_226 VSS VDD scs8hd_decap_4
XFILLER_16_12 VDD VSS scs8hd_fill_2
XFILLER_12_148 VSS VDD scs8hd_fill_1
XFILLER_16_78 VSS VDD scs8hd_decap_12
XANTENNA__515__A _515_/A VSS VDD scs8hd_diode_2
XFILLER_32_77 VSS VDD scs8hd_decap_8
X_675_ _667_/CLK _579_/X _574_/A _377_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__450__A1N _445_/Y VSS VDD scs8hd_diode_2
XANTENNA__425__A _366_/A VSS VDD scs8hd_diode_2
XFILLER_11_181 VDD VSS scs8hd_fill_2
XANTENNA__335__A _332_/X VSS VDD scs8hd_diode_2
XANTENNA__479__B2 _480_/B VSS VDD scs8hd_diode_2
X_391_ _389_/A _391_/X VSS VDD scs8hd_buf_1
XFILLER_27_55 VDD VSS scs8hd_fill_2
XFILLER_25_240 VSS VDD scs8hd_decap_4
X_460_ _460_/A _460_/Y VSS VDD scs8hd_inv_8
XFILLER_17_218 VDD VSS scs8hd_fill_2
XFILLER_40_232 VSS VDD scs8hd_fill_1
XFILLER_4_144 VSS VDD scs8hd_fill_1
XFILLER_4_48 VDD VSS scs8hd_fill_2
XFILLER_4_37 VDD VSS scs8hd_fill_2
XFILLER_4_26 VSS VDD scs8hd_decap_4
XFILLER_4_15 VSS VDD scs8hd_decap_4
XANTENNA__648__CLK _648_/CLK VSS VDD scs8hd_diode_2
X_589_ _682_/Q _589_/Y VSS VDD scs8hd_inv_8
XFILLER_31_243 VSS VDD scs8hd_fill_1
X_658_ _651_/CLK _515_/X _658_/Q _397_/X VSS VDD scs8hd_dfrtp_4
XFILLER_22_243 VSS VDD scs8hd_decap_8
XFILLER_1_103 VDD VSS scs8hd_fill_2
XFILLER_1_136 VDD VSS scs8hd_fill_2
XFILLER_38_98 VDD VSS scs8hd_fill_2
XFILLER_38_32 VSS VDD scs8hd_decap_3
XFILLER_38_21 VSS VDD scs8hd_decap_8
X_374_ _402_/A _375_/A VSS VDD scs8hd_buf_1
X_443_ _438_/Y _439_/Y _441_/X _442_/X _443_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_13_210 VDD VSS scs8hd_fill_2
X_512_ _512_/A _515_/A VSS VDD scs8hd_buf_1
XFILLER_0_180 VDD VSS scs8hd_fill_2
XANTENNA__645__RESETB _412_/X VSS VDD scs8hd_diode_2
XANTENNA__615__B2 _616_/B VSS VDD scs8hd_diode_2
XANTENNA__613__A _612_/X VSS VDD scs8hd_diode_2
XFILLER_39_184 VSS VDD scs8hd_decap_4
XANTENNA__542__B1 _538_/A VSS VDD scs8hd_diode_2
XFILLER_10_224 VSS VDD scs8hd_decap_4
XFILLER_10_235 VSS VDD scs8hd_decap_4
XANTENNA__523__A _520_/X VSS VDD scs8hd_diode_2
XFILLER_40_88 VSS VDD scs8hd_decap_4
XFILLER_6_3 VDD VSS scs8hd_fill_2
X_426_ _633_/Q _426_/Y VSS VDD scs8hd_inv_8
X_357_ _357_/A _357_/X VSS VDD scs8hd_buf_1
XANTENNA__486__A2N _482_/Y VSS VDD scs8hd_diode_2
XFILLER_39_3 VDD VSS scs8hd_fill_2
XFILLER_36_154 VSS VDD scs8hd_decap_3
XANTENNA__343__A _343_/A VSS VDD scs8hd_diode_2
XFILLER_19_12 VDD VSS scs8hd_fill_2
XFILLER_27_154 VDD VSS scs8hd_fill_2
XFILLER_19_34 VSS VDD scs8hd_fill_1
XFILLER_19_45 VSS VDD scs8hd_fill_1
XFILLER_42_146 VSS VDD scs8hd_decap_8
XFILLER_35_88 VDD VSS scs8hd_fill_2
XANTENNA__518__A _518_/A VSS VDD scs8hd_diode_2
XANTENNA__557__A1N _552_/Y VSS VDD scs8hd_diode_2
XANTENNA__428__A y VSS VDD scs8hd_diode_2
XFILLER_18_154 VDD VSS scs8hd_fill_2
X_409_ _402_/A _410_/A VSS VDD scs8hd_buf_1
XANTENNA__506__B1 _502_/A VSS VDD scs8hd_diode_2
XFILLER_24_102 VSS VDD scs8hd_decap_3
XFILLER_2_81 VDD VSS scs8hd_fill_2
XPHY_108 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__338__A _605_/A VSS VDD scs8hd_diode_2
XPHY_119 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__681__CLK _681_/CLK VSS VDD scs8hd_diode_2
X_691_ _681_/CLK _691_/D _691_/Q _356_/X VSS VDD scs8hd_dfrtp_4
XFILLER_30_127 VDD VSS scs8hd_fill_2
XFILLER_7_37 VSS VDD scs8hd_decap_3
XFILLER_7_48 VDD VSS scs8hd_fill_2
XFILLER_7_59 VDD VSS scs8hd_fill_2
XFILLER_30_7 VDD VSS scs8hd_fill_2
XANTENNA__430__B x[0] VSS VDD scs8hd_diode_2
XFILLER_14_190 VDD VSS scs8hd_fill_2
XANTENNA__605__B x[24] VSS VDD scs8hd_diode_2
XANTENNA__693__RESETB _354_/X VSS VDD scs8hd_diode_2
XFILLER_16_24 VSS VDD scs8hd_decap_3
XFILLER_32_23 VDD VSS scs8hd_fill_2
XFILLER_32_12 VDD VSS scs8hd_fill_2
XANTENNA__515__B _513_/X VSS VDD scs8hd_diode_2
XFILLER_20_182 VDD VSS scs8hd_fill_2
XANTENNA__531__A _663_/Q VSS VDD scs8hd_diode_2
X_674_ _667_/CLK _674_/D _560_/A _378_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_142 VDD VSS scs8hd_fill_2
XFILLER_11_171 VSS VDD scs8hd_decap_4
XANTENNA__441__A _441_/A VSS VDD scs8hd_diode_2
XFILLER_21_3 VDD VSS scs8hd_fill_2
XFILLER_26_219 VSS VDD scs8hd_decap_4
XFILLER_26_208 VDD VSS scs8hd_fill_2
XANTENNA__335__B _333_/X VSS VDD scs8hd_diode_2
XANTENNA__616__A _616_/A VSS VDD scs8hd_diode_2
XANTENNA__351__A rst VSS VDD scs8hd_diode_2
XFILLER_8_91 VSS VDD scs8hd_fill_1
XFILLER_27_34 VDD VSS scs8hd_fill_2
X_390_ _389_/A _390_/X VSS VDD scs8hd_buf_1
XANTENNA__526__A _547_/A VSS VDD scs8hd_diode_2
XFILLER_4_123 VDD VSS scs8hd_fill_2
XFILLER_4_189 VDD VSS scs8hd_fill_2
XFILLER_16_241 VSS VDD scs8hd_decap_12
X_657_ _651_/CLK _514_/X _657_/Q _398_/X VSS VDD scs8hd_dfrtp_4
X_588_ _679_/Q _588_/Y VSS VDD scs8hd_inv_8
XFILLER_31_233 VDD VSS scs8hd_fill_2
XANTENNA__641__RESETB _417_/X VSS VDD scs8hd_diode_2
XANTENNA__436__A _635_/Q VSS VDD scs8hd_diode_2
XANTENNA__346__A _345_/X VSS VDD scs8hd_diode_2
XFILLER_13_47 VDD VSS scs8hd_fill_2
XFILLER_38_66 VSS VDD scs8hd_decap_4
X_511_ _476_/A x[11] _512_/A VSS VDD scs8hd_and2_4
X_442_ _438_/Y _439_/Y _438_/A _640_/Q _442_/X VSS VDD scs8hd_o22a_4
X_373_ _373_/A _402_/A VSS VDD scs8hd_buf_1
XFILLER_0_192 VDD VSS scs8hd_fill_2
XANTENNA__608__A2N _603_/Y VSS VDD scs8hd_diode_2
XFILLER_5_92 VSS VDD scs8hd_decap_4
XFILLER_24_68 VDD VSS scs8hd_fill_2
XFILLER_40_12 VSS VDD scs8hd_decap_3
XANTENNA__542__A1 _538_/Y VSS VDD scs8hd_diode_2
XANTENNA__542__B2 _539_/A VSS VDD scs8hd_diode_2
XANTENNA__638__CLK _648_/CLK VSS VDD scs8hd_diode_2
XANTENNA__523__B _521_/X VSS VDD scs8hd_diode_2
XFILLER_1_17 VSS VDD scs8hd_decap_4
XFILLER_1_39 VSS VDD scs8hd_decap_4
X_425_ _366_/A _425_/X VSS VDD scs8hd_buf_1
X_356_ _357_/A _356_/X VSS VDD scs8hd_buf_1
XANTENNA__486__A1N _481_/Y VSS VDD scs8hd_diode_2
XFILLER_36_111 VDD VSS scs8hd_fill_2
XFILLER_36_177 VSS VDD scs8hd_fill_1
XFILLER_10_26 VSS VDD scs8hd_decap_4
XFILLER_10_37 VSS VDD scs8hd_decap_6
XANTENNA__624__A _624_/A VSS VDD scs8hd_diode_2
XFILLER_19_24 VDD VSS scs8hd_fill_2
XFILLER_42_125 VSS VDD scs8hd_decap_4
XFILLER_35_34 VDD VSS scs8hd_fill_2
XFILLER_35_23 VDD VSS scs8hd_fill_2
XFILLER_27_177 VDD VSS scs8hd_fill_2
XFILLER_27_111 VDD VSS scs8hd_fill_2
XANTENNA__534__A _533_/X VSS VDD scs8hd_diode_2
XANTENNA__688__RESETB _361_/X VSS VDD scs8hd_diode_2
XFILLER_2_210 VSS VDD scs8hd_decap_4
X_408_ _405_/A _408_/X VSS VDD scs8hd_buf_1
XFILLER_18_199 VSS VDD scs8hd_decap_4
XANTENNA__506__A1 _502_/Y VSS VDD scs8hd_diode_2
XANTENNA__444__A _441_/X VSS VDD scs8hd_diode_2
X_339_ _339_/A _339_/X VSS VDD scs8hd_buf_1
XANTENNA__506__B2 _658_/Q VSS VDD scs8hd_diode_2
XFILLER_24_125 VSS VDD scs8hd_decap_3
XFILLER_2_93 VSS VDD scs8hd_decap_6
XANTENNA__619__A _605_/A VSS VDD scs8hd_diode_2
XANTENNA__338__B x[29] VSS VDD scs8hd_diode_2
XANTENNA__442__B1 _438_/A VSS VDD scs8hd_diode_2
XFILLER_24_169 VDD VSS scs8hd_fill_2
XFILLER_24_147 VSS VDD scs8hd_decap_6
XPHY_109 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__354__A _357_/A VSS VDD scs8hd_diode_2
X_690_ _681_/CLK _630_/X _690_/Q _357_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__433__B1 _434_/A VSS VDD scs8hd_diode_2
XFILLER_15_114 VDD VSS scs8hd_fill_2
XFILLER_15_136 VSS VDD scs8hd_decap_4
XFILLER_23_7 VSS VDD scs8hd_fill_1
XFILLER_11_91 VDD VSS scs8hd_fill_2
XFILLER_38_206 VSS VDD scs8hd_decap_8
XANTENNA__439__A _640_/Q VSS VDD scs8hd_diode_2
XFILLER_21_106 VDD VSS scs8hd_fill_2
XANTENNA__636__RESETB _422_/X VSS VDD scs8hd_diode_2
XANTENNA__349__A _346_/X VSS VDD scs8hd_diode_2
XFILLER_16_36 VSS VDD scs8hd_decap_3
XFILLER_32_46 VSS VDD scs8hd_decap_4
XFILLER_20_172 VDD VSS scs8hd_fill_2
XFILLER_35_209 VDD VSS scs8hd_fill_2
X_673_ _667_/CLK _572_/X _673_/Q _379_/X VSS VDD scs8hd_dfrtp_4
XFILLER_22_90 VDD VSS scs8hd_fill_2
XFILLER_14_3 VSS VDD scs8hd_decap_4
XFILLER_34_220 VDD VSS scs8hd_fill_2
XANTENNA__632__A _694_/Q VSS VDD scs8hd_diode_2
XANTENNA__616__B _616_/B VSS VDD scs8hd_diode_2
XANTENNA__671__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_17_209 VDD VSS scs8hd_fill_2
XFILLER_27_79 VSS VDD scs8hd_fill_1
XANTENNA__526__B x[13] VSS VDD scs8hd_diode_2
XANTENNA__514__A2N _510_/Y VSS VDD scs8hd_diode_2
XFILLER_4_179 VSS VDD scs8hd_decap_3
X_587_ _584_/X _587_/B _587_/X VSS VDD scs8hd_xor2_4
X_656_ _651_/CLK _508_/X _496_/A _399_/X VSS VDD scs8hd_dfrtp_4
XFILLER_16_220 VDD VSS scs8hd_fill_2
XFILLER_17_90 VDD VSS scs8hd_fill_2
XFILLER_31_245 VSS VDD scs8hd_decap_8
XANTENNA__436__B _435_/X VSS VDD scs8hd_diode_2
XANTENNA__694__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__452__A _452_/A VSS VDD scs8hd_diode_2
XFILLER_22_212 VDD VSS scs8hd_fill_2
XANTENNA__627__A _626_/X VSS VDD scs8hd_diode_2
XFILLER_13_15 VDD VSS scs8hd_fill_2
XANTENNA__362__A _363_/A VSS VDD scs8hd_diode_2
XFILLER_13_59 VDD VSS scs8hd_fill_2
XANTENNA__537__A _534_/X VSS VDD scs8hd_diode_2
X_441_ _441_/A _441_/X VSS VDD scs8hd_buf_1
X_510_ _660_/Q _510_/Y VSS VDD scs8hd_inv_8
X_372_ _370_/A _372_/X VSS VDD scs8hd_buf_1
XFILLER_13_245 VDD VSS scs8hd_fill_2
X_639_ _648_/CLK _450_/X _445_/A _419_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__447__A _461_/A VSS VDD scs8hd_diode_2
XANTENNA__608__A1N _602_/Y VSS VDD scs8hd_diode_2
XFILLER_39_120 VDD VSS scs8hd_fill_2
XANTENNA__357__A _357_/A VSS VDD scs8hd_diode_2
XFILLER_24_36 VDD VSS scs8hd_fill_2
XFILLER_24_25 VDD VSS scs8hd_fill_2
XFILLER_10_215 VDD VSS scs8hd_fill_2
XANTENNA__542__A2 _539_/Y VSS VDD scs8hd_diode_2
XANTENNA__684__RESETB _365_/X VSS VDD scs8hd_diode_2
X_424_ _366_/A _424_/X VSS VDD scs8hd_buf_1
X_355_ _357_/A _355_/X VSS VDD scs8hd_buf_1
XFILLER_14_91 VSS VDD scs8hd_fill_1
XFILLER_30_90 VDD VSS scs8hd_fill_2
XFILLER_36_167 VSS VDD scs8hd_fill_1
XFILLER_36_145 VDD VSS scs8hd_fill_2
XFILLER_36_134 VDD VSS scs8hd_fill_2
XFILLER_42_104 VSS VDD scs8hd_fill_1
XFILLER_35_46 VSS VDD scs8hd_decap_12
XFILLER_27_134 VSS VDD scs8hd_decap_4
XFILLER_27_123 VSS VDD scs8hd_decap_4
XFILLER_18_123 VDD VSS scs8hd_fill_2
XFILLER_18_134 VDD VSS scs8hd_fill_2
XFILLER_18_167 VSS VDD scs8hd_decap_12
XFILLER_41_181 VDD VSS scs8hd_fill_2
X_407_ _405_/A _407_/X VSS VDD scs8hd_buf_1
XANTENNA__444__B _442_/X VSS VDD scs8hd_diode_2
XPHY_90 VSS VDD scs8hd_tapvpwrvgnd_1
X_338_ _605_/A x[29] _339_/A VSS VDD scs8hd_and2_4
XANTENNA__460__A _460_/A VSS VDD scs8hd_diode_2
XANTENNA__506__A2 _503_/Y VSS VDD scs8hd_diode_2
XFILLER_24_137 VSS VDD scs8hd_decap_8
XANTENNA__619__B x[26] VSS VDD scs8hd_diode_2
XANTENNA__442__B2 _640_/Q VSS VDD scs8hd_diode_2
XANTENNA__442__A1 _438_/Y VSS VDD scs8hd_diode_2
XFILLER_21_15 VDD VSS scs8hd_fill_2
XANTENNA__370__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_21_59 VDD VSS scs8hd_fill_2
XANTENNA__433__B2 _434_/B VSS VDD scs8hd_diode_2
XANTENNA__545__A _545_/A VSS VDD scs8hd_diode_2
XFILLER_23_181 VDD VSS scs8hd_fill_2
XFILLER_14_170 VDD VSS scs8hd_fill_2
XANTENNA__455__A _454_/X VSS VDD scs8hd_diode_2
XFILLER_37_240 VSS VDD scs8hd_decap_4
XANTENNA__349__B _347_/X VSS VDD scs8hd_diode_2
XANTENNA__365__A _363_/A VSS VDD scs8hd_diode_2
XFILLER_32_36 VSS VDD scs8hd_fill_1
XFILLER_20_151 VDD VSS scs8hd_fill_2
XANTENNA__443__A2N _439_/Y VSS VDD scs8hd_diode_2
XANTENNA__593__A2N _589_/Y VSS VDD scs8hd_diode_2
X_672_ _667_/CLK _672_/D _553_/A _380_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_177 VDD VSS scs8hd_fill_2
XFILLER_11_184 VDD VSS scs8hd_fill_2
XANTENNA__333__B1 _691_/Q VSS VDD scs8hd_diode_2
XFILLER_8_93 VDD VSS scs8hd_fill_2
XFILLER_25_221 VDD VSS scs8hd_fill_2
XANTENNA__572__B1 _570_/X VSS VDD scs8hd_diode_2
XANTENNA__514__A1N _509_/Y VSS VDD scs8hd_diode_2
XFILLER_4_147 VDD VSS scs8hd_fill_2
XFILLER_4_136 VSS VDD scs8hd_decap_8
XFILLER_4_114 VSS VDD scs8hd_decap_6
X_586_ _581_/Y _582_/Y _584_/X _587_/B _586_/X VSS VDD scs8hd_a2bb2o_4
X_655_ _651_/CLK _507_/X _502_/A _400_/X VSS VDD scs8hd_dfrtp_4
XPHY_260 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__679__RESETB _371_/X VSS VDD scs8hd_diode_2
XFILLER_38_13 VDD VSS scs8hd_fill_2
XFILLER_1_117 VSS VDD scs8hd_fill_1
XANTENNA__537__B _535_/X VSS VDD scs8hd_diode_2
X_371_ _370_/A _371_/X VSS VDD scs8hd_buf_1
X_440_ _461_/A x[1] _441_/A VSS VDD scs8hd_and2_4
XFILLER_13_224 VSS VDD scs8hd_fill_1
XANTENNA__680__RESETB _370_/X VSS VDD scs8hd_diode_2
XANTENNA__553__A _553_/A VSS VDD scs8hd_diode_2
XFILLER_28_90 VDD VSS scs8hd_fill_2
XFILLER_0_150 VSS VDD scs8hd_decap_4
XANTENNA__536__B1 _534_/X VSS VDD scs8hd_diode_2
XANTENNA__661__CLK _651_/CLK VSS VDD scs8hd_diode_2
X_638_ _648_/CLK _444_/X _638_/Q _420_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__447__B x[2] VSS VDD scs8hd_diode_2
X_569_ _597_/A x[19] _570_/A VSS VDD scs8hd_and2_4
XFILLER_39_176 VDD VSS scs8hd_fill_2
XFILLER_39_154 VDD VSS scs8hd_fill_2
XFILLER_6_209 VSS VDD scs8hd_fill_1
XANTENNA__373__A _373_/A VSS VDD scs8hd_diode_2
XFILLER_40_58 VDD VSS scs8hd_fill_2
XFILLER_40_69 VDD VSS scs8hd_fill_2
XANTENNA__548__A _547_/X VSS VDD scs8hd_diode_2
XANTENNA__684__CLK _681_/CLK VSS VDD scs8hd_diode_2
X_354_ _357_/A _354_/X VSS VDD scs8hd_buf_1
X_423_ _366_/A _423_/X VSS VDD scs8hd_buf_1
XFILLER_14_70 VDD VSS scs8hd_fill_2
XFILLER_14_81 VDD VSS scs8hd_fill_2
XANTENNA__458__A _458_/A VSS VDD scs8hd_diode_2
XANTENNA__368__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_19_37 VDD VSS scs8hd_fill_2
XFILLER_19_59 VDD VSS scs8hd_fill_2
XFILLER_42_138 VDD VSS scs8hd_fill_2
XFILLER_35_58 VSS VDD scs8hd_decap_3
XFILLER_4_3 VDD VSS scs8hd_fill_2
XFILLER_2_201 VDD VSS scs8hd_fill_2
XFILLER_33_127 VSS VDD scs8hd_decap_4
XFILLER_18_146 VSS VDD scs8hd_decap_3
XFILLER_18_179 VSS VDD scs8hd_fill_1
XFILLER_41_171 VSS VDD scs8hd_decap_4
XPHY_80 VSS VDD scs8hd_decap_3
XFILLER_33_138 VDD VSS scs8hd_fill_2
X_406_ _405_/A _406_/X VSS VDD scs8hd_buf_1
XPHY_91 VSS VDD scs8hd_tapvpwrvgnd_1
X_337_ _337_/A _337_/Y VSS VDD scs8hd_inv_8
XFILLER_37_3 VSS VDD scs8hd_decap_4
XFILLER_2_51 VDD VSS scs8hd_fill_2
XANTENNA__442__A2 _439_/Y VSS VDD scs8hd_diode_2
XFILLER_32_171 VDD VSS scs8hd_fill_2
XANTENNA__561__A _518_/A VSS VDD scs8hd_diode_2
XFILLER_38_219 VSS VDD scs8hd_fill_1
XFILLER_16_8 VDD VSS scs8hd_fill_2
XFILLER_36_90 VDD VSS scs8hd_fill_2
XFILLER_16_16 VDD VSS scs8hd_fill_2
XFILLER_20_141 VSS VDD scs8hd_fill_1
XANTENNA__381__A _402_/A VSS VDD scs8hd_diode_2
XANTENNA__443__A1N _438_/Y VSS VDD scs8hd_diode_2
XANTENNA__593__A1N _588_/Y VSS VDD scs8hd_diode_2
XFILLER_28_252 VSS VDD scs8hd_fill_1
X_671_ _667_/CLK _565_/X _671_/Q _382_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_123 VDD VSS scs8hd_fill_2
XFILLER_11_141 VDD VSS scs8hd_fill_2
XFILLER_11_152 VSS VDD scs8hd_decap_3
XFILLER_11_163 VDD VSS scs8hd_fill_2
XANTENNA__675__RESETB _377_/X VSS VDD scs8hd_diode_2
XANTENNA__466__A _645_/Q VSS VDD scs8hd_diode_2
XANTENNA__333__B2 _694_/Q VSS VDD scs8hd_diode_2
XANTENNA__333__A1 _631_/Y VSS VDD scs8hd_diode_2
XFILLER_27_59 VDD VSS scs8hd_fill_2
XANTENNA__376__A _375_/A VSS VDD scs8hd_diode_2
XANTENNA__572__B2 _573_/B VSS VDD scs8hd_diode_2
XFILLER_4_19 VSS VDD scs8hd_fill_1
X_654_ _651_/CLK _501_/X _489_/A _401_/X VSS VDD scs8hd_dfrtp_4
XPHY_261 VSS VDD scs8hd_tapvpwrvgnd_1
X_585_ _581_/Y _582_/Y _581_/A _582_/A _587_/B VSS VDD scs8hd_o22a_4
XPHY_250 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_31_225 VSS VDD scs8hd_fill_1
XFILLER_3_181 VDD VSS scs8hd_fill_2
XANTENNA__433__A2N _427_/Y VSS VDD scs8hd_diode_2
XFILLER_1_107 VSS VDD scs8hd_decap_3
X_370_ _370_/A _370_/X VSS VDD scs8hd_buf_1
XFILLER_9_207 VDD VSS scs8hd_fill_2
XFILLER_13_214 VDD VSS scs8hd_fill_2
XFILLER_13_236 VDD VSS scs8hd_fill_2
XFILLER_0_184 VDD VSS scs8hd_fill_2
X_637_ _648_/CLK _443_/X _438_/A _421_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__536__B2 _535_/X VSS VDD scs8hd_diode_2
X_499_ _495_/Y _496_/Y _653_/Q _496_/A _501_/B VSS VDD scs8hd_o22a_4
X_568_ _676_/Q _568_/Y VSS VDD scs8hd_inv_8
XFILLER_5_62 VSS VDD scs8hd_decap_3
XFILLER_5_51 VDD VSS scs8hd_fill_2
XFILLER_10_206 VDD VSS scs8hd_fill_2
XFILLER_6_7 VDD VSS scs8hd_fill_2
XANTENNA__479__A2N _474_/Y VSS VDD scs8hd_diode_2
XANTENNA__463__B1 _643_/Q VSS VDD scs8hd_diode_2
X_353_ _357_/A _353_/X VSS VDD scs8hd_buf_1
X_422_ _417_/A _422_/X VSS VDD scs8hd_buf_1
XFILLER_5_243 VSS VDD scs8hd_fill_1
XFILLER_14_93 VDD VSS scs8hd_fill_2
XFILLER_39_7 VDD VSS scs8hd_fill_2
XANTENNA__474__A _474_/A VSS VDD scs8hd_diode_2
XANTENNA__458__B _456_/X VSS VDD scs8hd_diode_2
XFILLER_27_158 VSS VDD scs8hd_decap_4
XFILLER_19_16 VDD VSS scs8hd_fill_2
XFILLER_19_49 VDD VSS scs8hd_fill_2
XANTENNA__384__A _386_/A VSS VDD scs8hd_diode_2
XANTENNA__651__CLK _651_/CLK VSS VDD scs8hd_diode_2
XANTENNA__559__A _671_/Q VSS VDD scs8hd_diode_2
XFILLER_18_158 VDD VSS scs8hd_fill_2
XFILLER_41_161 VDD VSS scs8hd_fill_2
XPHY_81 VSS VDD scs8hd_decap_3
X_405_ _405_/A _405_/X VSS VDD scs8hd_buf_1
XPHY_70 VSS VDD scs8hd_decap_3
X_336_ _693_/Q _336_/Y VSS VDD scs8hd_inv_8
XPHY_92 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__469__A _469_/A VSS VDD scs8hd_diode_2
XFILLER_2_85 VSS VDD scs8hd_decap_6
XANTENNA__674__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__379__A _375_/A VSS VDD scs8hd_diode_2
XFILLER_15_106 VDD VSS scs8hd_fill_2
XFILLER_15_128 VDD VSS scs8hd_fill_2
XANTENNA__671__RESETB _382_/X VSS VDD scs8hd_diode_2
XFILLER_14_194 VSS VDD scs8hd_decap_12
XFILLER_32_27 VSS VDD scs8hd_decap_4
XFILLER_12_109 VDD VSS scs8hd_fill_2
XFILLER_20_186 VDD VSS scs8hd_fill_2
XFILLER_20_197 VDD VSS scs8hd_fill_2
X_670_ _667_/CLK _670_/D _546_/A _383_/X VSS VDD scs8hd_dfrtp_4
XFILLER_22_93 VSS VDD scs8hd_decap_4
XFILLER_22_82 VSS VDD scs8hd_decap_8
XFILLER_7_146 VDD VSS scs8hd_fill_2
XFILLER_11_120 VDD VSS scs8hd_fill_2
XFILLER_34_212 VDD VSS scs8hd_fill_2
XANTENNA__482__A _652_/Q VSS VDD scs8hd_diode_2
XFILLER_34_245 VSS VDD scs8hd_decap_8
XANTENNA__333__A2 _632_/Y VSS VDD scs8hd_diode_2
XFILLER_6_190 VSS VDD scs8hd_decap_4
XFILLER_8_62 VDD VSS scs8hd_fill_2
XFILLER_40_226 VSS VDD scs8hd_decap_6
XFILLER_40_215 VDD VSS scs8hd_fill_2
XFILLER_27_38 VSS VDD scs8hd_decap_4
XFILLER_25_245 VSS VDD scs8hd_decap_8
XANTENNA__392__A _389_/A VSS VDD scs8hd_diode_2
XFILLER_4_127 VDD VSS scs8hd_fill_2
X_653_ _651_/CLK _653_/D _653_/Q _403_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__567__A _673_/Q VSS VDD scs8hd_diode_2
XFILLER_16_212 VDD VSS scs8hd_fill_2
XPHY_262 VSS VDD scs8hd_tapvpwrvgnd_1
X_584_ _583_/X _584_/X VSS VDD scs8hd_buf_1
XPHY_251 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_240 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_31_237 VSS VDD scs8hd_decap_6
XFILLER_12_3 VDD VSS scs8hd_fill_2
XANTENNA__477__A _476_/X VSS VDD scs8hd_diode_2
XFILLER_22_215 VSS VDD scs8hd_decap_4
XANTENNA__433__A1N _426_/Y VSS VDD scs8hd_diode_2
XFILLER_38_37 VDD VSS scs8hd_fill_2
XANTENNA__387__A _386_/A VSS VDD scs8hd_diode_2
XFILLER_13_204 VSS VDD scs8hd_decap_3
XFILLER_0_196 VSS VDD scs8hd_decap_4
XFILLER_0_130 VDD VSS scs8hd_fill_2
X_636_ _648_/CLK _437_/Y _344_/A _422_/X VSS VDD scs8hd_dfrtp_4
X_567_ _673_/Q _567_/Y VSS VDD scs8hd_inv_8
X_498_ _497_/X _498_/X VSS VDD scs8hd_buf_1
XFILLER_39_123 VDD VSS scs8hd_fill_2
XFILLER_39_112 VDD VSS scs8hd_fill_2
XANTENNA__550__A2N _546_/Y VSS VDD scs8hd_diode_2
XANTENNA__479__A1N _473_/Y VSS VDD scs8hd_diode_2
X_421_ _417_/A _421_/X VSS VDD scs8hd_buf_1
XANTENNA__463__A1 _459_/Y VSS VDD scs8hd_diode_2
XANTENNA__463__B2 _460_/A VSS VDD scs8hd_diode_2
X_352_ _373_/A _357_/A VSS VDD scs8hd_buf_1
XFILLER_30_93 VSS VDD scs8hd_decap_3
XFILLER_5_222 VDD VSS scs8hd_fill_2
XFILLER_5_233 VDD VSS scs8hd_fill_2
XANTENNA__580__A _580_/A VSS VDD scs8hd_diode_2
XFILLER_36_126 VDD VSS scs8hd_fill_2
XFILLER_36_115 VDD VSS scs8hd_fill_2
XFILLER_36_159 VDD VSS scs8hd_fill_2
X_619_ _605_/A x[26] _620_/A VSS VDD scs8hd_and2_4
XANTENNA__490__A _476_/A VSS VDD scs8hd_diode_2
XANTENNA__666__RESETB _387_/X VSS VDD scs8hd_diode_2
XANTENNA__640__D _451_/X VSS VDD scs8hd_diode_2
XFILLER_19_28 VSS VDD scs8hd_decap_6
XFILLER_42_107 VSS VDD scs8hd_decap_12
XFILLER_35_38 VDD VSS scs8hd_fill_2
XFILLER_35_27 VSS VDD scs8hd_decap_4
XFILLER_27_115 VSS VDD scs8hd_decap_3
XFILLER_35_181 VDD VSS scs8hd_fill_2
XFILLER_35_170 VSS VDD scs8hd_decap_4
XPHY_82 VSS VDD scs8hd_decap_3
XPHY_71 VSS VDD scs8hd_decap_3
X_404_ _405_/A _404_/X VSS VDD scs8hd_buf_1
XFILLER_33_107 VDD VSS scs8hd_fill_2
XPHY_60 VSS VDD scs8hd_decap_3
XFILLER_26_192 VSS VDD scs8hd_decap_3
XANTENNA__575__A _678_/Q VSS VDD scs8hd_diode_2
XFILLER_41_184 VDD VSS scs8hd_fill_2
XFILLER_25_93 VSS VDD scs8hd_fill_1
X_335_ _332_/X _333_/X _692_/D VSS VDD scs8hd_xor2_4
XPHY_93 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_24_107 VDD VSS scs8hd_fill_2
XFILLER_32_195 VDD VSS scs8hd_fill_2
XANTENNA__635__D _436_/X VSS VDD scs8hd_diode_2
XFILLER_17_181 VDD VSS scs8hd_fill_2
XANTENNA__395__A _402_/A VSS VDD scs8hd_diode_2
XFILLER_15_118 VSS VDD scs8hd_decap_4
XFILLER_23_184 VDD VSS scs8hd_fill_2
XFILLER_23_162 VSS VDD scs8hd_decap_4
XFILLER_11_62 VDD VSS scs8hd_fill_2
XANTENNA__593__B1 _594_/A VSS VDD scs8hd_diode_2
XFILLER_14_151 VDD VSS scs8hd_fill_2
XFILLER_42_3 VSS VDD scs8hd_decap_12
XFILLER_16_29 VDD VSS scs8hd_fill_2
XANTENNA__641__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_20_154 VDD VSS scs8hd_fill_2
XFILLER_20_176 VSS VDD scs8hd_decap_4
XFILLER_11_132 VSS VDD scs8hd_decap_6
XFILLER_22_61 VDD VSS scs8hd_fill_2
XFILLER_22_50 VSS VDD scs8hd_decap_4
XFILLER_7_103 VSS VDD scs8hd_decap_4
XFILLER_7_114 VDD VSS scs8hd_fill_2
XFILLER_21_8 VSS VDD scs8hd_decap_4
XANTENNA__664__CLK _651_/CLK VSS VDD scs8hd_diode_2
XANTENNA__507__A2N _503_/Y VSS VDD scs8hd_diode_2
XANTENNA__557__B1 _558_/A VSS VDD scs8hd_diode_2
XFILLER_25_213 VDD VSS scs8hd_fill_2
X_583_ _597_/A x[21] _583_/X VSS VDD scs8hd_and2_4
X_652_ _651_/CLK _494_/X _652_/Q _404_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__687__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_16_224 VSS VDD scs8hd_decap_3
XFILLER_17_50 VSS VDD scs8hd_decap_8
XFILLER_17_72 VSS VDD scs8hd_fill_1
XPHY_263 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__583__A _597_/A VSS VDD scs8hd_diode_2
XPHY_252 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_241 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_230 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_71 VDD VSS scs8hd_fill_2
XFILLER_33_60 VSS VDD scs8hd_fill_1
XFILLER_3_172 VDD VSS scs8hd_fill_2
XANTENNA__643__D _643_/D VSS VDD scs8hd_diode_2
XFILLER_13_227 VDD VSS scs8hd_fill_2
XFILLER_13_249 VSS VDD scs8hd_decap_4
XFILLER_0_142 VDD VSS scs8hd_fill_2
XFILLER_28_93 VDD VSS scs8hd_fill_2
X_566_ _566_/A _566_/B _672_/D VSS VDD scs8hd_xor2_4
X_635_ _648_/CLK _436_/X _635_/Q _423_/X VSS VDD scs8hd_dfrtp_4
X_497_ _476_/A x[9] _497_/X VSS VDD scs8hd_and2_4
XFILLER_8_220 VDD VSS scs8hd_fill_2
XFILLER_5_42 VSS VDD scs8hd_decap_3
XFILLER_5_31 VSS VDD scs8hd_fill_1
XANTENNA__488__A _488_/A VSS VDD scs8hd_diode_2
XANTENNA__638__D _444_/X VSS VDD scs8hd_diode_2
XANTENNA__550__A1N _545_/Y VSS VDD scs8hd_diode_2
XANTENNA__662__RESETB _392_/X VSS VDD scs8hd_diode_2
XFILLER_24_29 VDD VSS scs8hd_fill_2
XFILLER_40_17 VSS VDD scs8hd_decap_12
XANTENNA__398__A _401_/A VSS VDD scs8hd_diode_2
XANTENNA__463__A2 _460_/Y VSS VDD scs8hd_diode_2
XFILLER_38_190 VDD VSS scs8hd_fill_2
X_420_ _417_/A _420_/X VSS VDD scs8hd_buf_1
X_351_ rst _373_/A VSS VDD scs8hd_inv_8
XFILLER_14_51 VSS VDD scs8hd_decap_3
XANTENNA__580__B _578_/X VSS VDD scs8hd_diode_2
XFILLER_5_245 VSS VDD scs8hd_decap_8
XFILLER_36_149 VSS VDD scs8hd_decap_4
XFILLER_36_138 VSS VDD scs8hd_decap_4
X_549_ _545_/Y _546_/Y _545_/A _546_/A _551_/B VSS VDD scs8hd_o22a_4
X_618_ _690_/Q _618_/Y VSS VDD scs8hd_inv_8
XANTENNA__490__B x[8] VSS VDD scs8hd_diode_2
XFILLER_42_119 VSS VDD scs8hd_fill_1
XFILLER_35_160 VSS VDD scs8hd_decap_3
XFILLER_2_215 VDD VSS scs8hd_fill_2
XFILLER_18_127 VSS VDD scs8hd_decap_4
XFILLER_18_138 VDD VSS scs8hd_fill_2
XPHY_83 VSS VDD scs8hd_decap_3
XPHY_72 VSS VDD scs8hd_decap_3
XFILLER_33_119 VSS VDD scs8hd_decap_3
XPHY_61 VSS VDD scs8hd_decap_3
X_403_ _405_/A _403_/X VSS VDD scs8hd_buf_1
XPHY_50 VSS VDD scs8hd_decap_3
X_334_ _631_/Y _632_/Y _332_/X _333_/X _691_/D VSS VDD scs8hd_a2bb2o_4
XPHY_94 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_41_82 VDD VSS scs8hd_fill_2
XANTENNA__591__A _590_/X VSS VDD scs8hd_diode_2
XFILLER_2_32 VSS VDD scs8hd_decap_4
XFILLER_32_163 VSS VDD scs8hd_decap_6
XFILLER_32_152 VSS VDD scs8hd_fill_1
XANTENNA__651__D _493_/X VSS VDD scs8hd_diode_2
XFILLER_2_3 VSS VDD scs8hd_decap_12
XFILLER_11_52 VSS VDD scs8hd_decap_4
XFILLER_36_71 VDD VSS scs8hd_fill_2
XFILLER_36_93 VDD VSS scs8hd_fill_2
XANTENNA__593__B2 _592_/X VSS VDD scs8hd_diode_2
XFILLER_14_163 VSS VDD scs8hd_decap_4
XFILLER_14_174 VDD VSS scs8hd_fill_2
XFILLER_37_211 VSS VDD scs8hd_decap_4
XFILLER_35_3 VDD VSS scs8hd_fill_2
XANTENNA__496__A _496_/A VSS VDD scs8hd_diode_2
XANTENNA__646__D _472_/X VSS VDD scs8hd_diode_2
XANTENNA__586__A2N _582_/Y VSS VDD scs8hd_diode_2
XFILLER_20_122 VSS VDD scs8hd_fill_1
XFILLER_20_133 VSS VDD scs8hd_decap_8
XFILLER_20_144 VSS VDD scs8hd_decap_4
XFILLER_28_244 VSS VDD scs8hd_decap_8
XFILLER_11_177 VDD VSS scs8hd_fill_2
XFILLER_34_203 VDD VSS scs8hd_fill_2
XFILLER_8_97 VDD VSS scs8hd_fill_2
XANTENNA__507__A1N _502_/Y VSS VDD scs8hd_diode_2
XFILLER_6_170 VDD VSS scs8hd_fill_2
XFILLER_40_206 VSS VDD scs8hd_decap_8
XANTENNA__557__B2 _558_/B VSS VDD scs8hd_diode_2
XFILLER_25_236 VDD VSS scs8hd_fill_2
XFILLER_25_225 VDD VSS scs8hd_fill_2
XANTENNA__493__B1 _491_/X VSS VDD scs8hd_diode_2
XANTENNA__CTS_buf_1_0_A _CTS_root/X VSS VDD scs8hd_diode_2
XANTENNA__657__RESETB _398_/X VSS VDD scs8hd_diode_2
X_582_ _582_/A _582_/Y VSS VDD scs8hd_inv_8
X_651_ _651_/CLK _493_/X _488_/A _405_/X VSS VDD scs8hd_dfrtp_4
XFILLER_31_217 VSS VDD scs8hd_decap_8
XFILLER_17_62 VDD VSS scs8hd_fill_2
XFILLER_17_84 VSS VDD scs8hd_decap_4
XPHY_264 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__583__B x[21] VSS VDD scs8hd_diode_2
XPHY_253 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_242 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_231 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_220 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_3_184 VDD VSS scs8hd_fill_2
XFILLER_22_206 VSS VDD scs8hd_decap_4
XFILLER_38_17 VDD VSS scs8hd_fill_2
XANTENNA__654__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_28_83 VSS VDD scs8hd_decap_4
XFILLER_28_72 VDD VSS scs8hd_fill_2
X_634_ _648_/CLK _634_/D p _424_/X VSS VDD scs8hd_dfrtp_4
XFILLER_0_187 VDD VSS scs8hd_fill_2
XFILLER_0_154 VSS VDD scs8hd_fill_1
XANTENNA__594__A _594_/A VSS VDD scs8hd_diode_2
X_496_ _496_/A _496_/Y VSS VDD scs8hd_inv_8
X_565_ _559_/Y _560_/Y _566_/A _566_/B _565_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_39_103 VDD VSS scs8hd_fill_2
XFILLER_5_98 VSS VDD scs8hd_decap_8
XANTENNA__457__B1 _458_/A VSS VDD scs8hd_diode_2
XANTENNA__654__D _501_/X VSS VDD scs8hd_diode_2
XFILLER_40_29 VDD VSS scs8hd_fill_2
XANTENNA__677__CLK _667_/CLK VSS VDD scs8hd_diode_2
X_350_ _366_/A _350_/X VSS VDD scs8hd_buf_1
XFILLER_14_74 VSS VDD scs8hd_decap_4
XFILLER_14_85 VSS VDD scs8hd_decap_6
XANTENNA__589__A _682_/Q VSS VDD scs8hd_diode_2
XFILLER_30_73 VSS VDD scs8hd_decap_12
XFILLER_30_62 VDD VSS scs8hd_fill_2
XFILLER_39_82 VDD VSS scs8hd_fill_2
XFILLER_29_180 VSS VDD scs8hd_decap_3
X_617_ _687_/Q _617_/Y VSS VDD scs8hd_inv_8
X_548_ _547_/X _548_/X VSS VDD scs8hd_buf_1
X_479_ _473_/Y _474_/Y _477_/X _480_/B _479_/X VSS VDD scs8hd_a2bb2o_4
XANTENNA__649__D _486_/X VSS VDD scs8hd_diode_2
XFILLER_4_7 VDD VSS scs8hd_fill_2
XPHY_84 VSS VDD scs8hd_decap_3
XFILLER_41_120 VDD VSS scs8hd_fill_2
XPHY_73 VSS VDD scs8hd_decap_3
XPHY_62 VSS VDD scs8hd_decap_3
X_402_ _402_/A _405_/A VSS VDD scs8hd_buf_1
XPHY_51 VSS VDD scs8hd_decap_3
XFILLER_25_62 VSS VDD scs8hd_decap_4
X_333_ _631_/Y _632_/Y _691_/Q _694_/Q _333_/X VSS VDD scs8hd_o22a_4
XPHY_95 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_40 VSS VDD scs8hd_decap_3
XFILLER_2_55 VSS VDD scs8hd_decap_4
XFILLER_2_22 VSS VDD scs8hd_decap_4
XFILLER_32_131 VSS VDD scs8hd_decap_8
XFILLER_32_120 VSS VDD scs8hd_decap_8
XFILLER_32_142 VDD VSS scs8hd_fill_2
XFILLER_23_175 VSS VDD scs8hd_decap_4
XFILLER_23_120 VDD VSS scs8hd_fill_2
XFILLER_11_20 VSS VDD scs8hd_fill_1
XFILLER_36_83 VSS VDD scs8hd_decap_4
XFILLER_36_61 VSS VDD scs8hd_decap_8
XFILLER_37_245 VSS VDD scs8hd_decap_8
XFILLER_28_3 VDD VSS scs8hd_fill_2
XANTENNA__586__A1N _581_/Y VSS VDD scs8hd_diode_2
XANTENNA__662__D _662_/D VSS VDD scs8hd_diode_2
XFILLER_28_212 VDD VSS scs8hd_fill_2
XANTENNA__653__RESETB _403_/X VSS VDD scs8hd_diode_2
XFILLER_7_127 VSS VDD scs8hd_decap_12
XFILLER_11_123 VDD VSS scs8hd_fill_2
XFILLER_11_167 VDD VSS scs8hd_fill_2
XANTENNA__597__A _597_/A VSS VDD scs8hd_diode_2
XFILLER_19_245 VSS VDD scs8hd_decap_8
XFILLER_34_215 VSS VDD scs8hd_decap_3
XFILLER_8_21 VDD VSS scs8hd_fill_2
XFILLER_8_32 VSS VDD scs8hd_decap_4
XFILLER_6_182 VDD VSS scs8hd_fill_2
XANTENNA__657__D _514_/X VSS VDD scs8hd_diode_2
XANTENNA__493__B2 _492_/X VSS VDD scs8hd_diode_2
X_650_ _651_/CLK _487_/X _474_/A _406_/X VSS VDD scs8hd_dfrtp_4
X_581_ _581_/A _581_/Y VSS VDD scs8hd_inv_8
XPHY_243 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_232 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_221 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_31_229 VDD VSS scs8hd_fill_2
XPHY_210 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_16_204 VDD VSS scs8hd_fill_2
XFILLER_16_215 VDD VSS scs8hd_fill_2
XPHY_265 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_254 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_62 VSS VDD scs8hd_decap_3
XFILLER_30_240 VSS VDD scs8hd_decap_12
XFILLER_38_29 VDD VSS scs8hd_fill_2
XFILLER_13_218 VSS VDD scs8hd_decap_6
XFILLER_0_122 VDD VSS scs8hd_fill_2
X_633_ _648_/CLK _633_/D _633_/Q _425_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__594__B _592_/X VSS VDD scs8hd_diode_2
X_495_ _653_/Q _495_/Y VSS VDD scs8hd_inv_8
X_564_ _559_/Y _560_/Y _671_/Q _560_/A _566_/B VSS VDD scs8hd_o22a_4
XFILLER_5_55 VDD VSS scs8hd_fill_2
XFILLER_39_148 VSS VDD scs8hd_decap_4
XFILLER_10_3 VDD VSS scs8hd_fill_2
XANTENNA__457__B2 _456_/X VSS VDD scs8hd_diode_2
XANTENNA__670__D _670_/D VSS VDD scs8hd_diode_2
XFILLER_30_41 VSS VDD scs8hd_decap_4
XFILLER_14_97 VDD VSS scs8hd_fill_2
XFILLER_30_85 VSS VDD scs8hd_decap_3
X_547_ _547_/A x[16] _547_/X VSS VDD scs8hd_and2_4
X_616_ _616_/A _616_/B _686_/D VSS VDD scs8hd_xor2_4
X_478_ _473_/Y _474_/Y _473_/A _474_/A _480_/B VSS VDD scs8hd_o22a_4
XANTENNA__665__D _543_/X VSS VDD scs8hd_diode_2
XFILLER_35_184 VDD VSS scs8hd_fill_2
XANTENNA__644__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_2_206 VDD VSS scs8hd_fill_2
X_401_ _401_/A _401_/X VSS VDD scs8hd_buf_1
XFILLER_26_151 VDD VSS scs8hd_fill_2
XFILLER_26_140 VDD VSS scs8hd_fill_2
XPHY_30 VSS VDD scs8hd_decap_3
XPHY_85 VSS VDD scs8hd_decap_3
XFILLER_41_165 VSS VDD scs8hd_decap_4
XFILLER_41_132 VDD VSS scs8hd_fill_2
XPHY_74 VSS VDD scs8hd_decap_3
XPHY_63 VSS VDD scs8hd_decap_3
XFILLER_26_184 VDD VSS scs8hd_fill_2
XPHY_52 VSS VDD scs8hd_decap_3
XFILLER_25_96 VDD VSS scs8hd_fill_2
XPHY_96 VSS VDD scs8hd_tapvpwrvgnd_1
X_332_ _331_/X _332_/X VSS VDD scs8hd_buf_1
XPHY_41 VSS VDD scs8hd_decap_3
XFILLER_41_73 VDD VSS scs8hd_fill_2
XFILLER_41_62 VSS VDD scs8hd_decap_4
XANTENNA__667__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__648__RESETB _408_/X VSS VDD scs8hd_diode_2
XFILLER_32_154 VDD VSS scs8hd_fill_2
XFILLER_32_110 VSS VDD scs8hd_fill_1
XFILLER_17_184 VDD VSS scs8hd_fill_2
XANTENNA__348__B1 _346_/X VSS VDD scs8hd_diode_2
XFILLER_23_154 VDD VSS scs8hd_fill_2
XFILLER_23_143 VDD VSS scs8hd_fill_2
XFILLER_11_87 VDD VSS scs8hd_fill_2
XFILLER_14_121 VDD VSS scs8hd_fill_2
XFILLER_14_154 VDD VSS scs8hd_fill_2
XANTENNA__578__B1 _574_/A VSS VDD scs8hd_diode_2
XFILLER_7_139 VSS VDD scs8hd_fill_1
XFILLER_11_113 VSS VDD scs8hd_decap_4
XFILLER_11_157 VSS VDD scs8hd_decap_3
XANTENNA__597__B x[23] VSS VDD scs8hd_diode_2
XFILLER_6_150 VSS VDD scs8hd_decap_3
XFILLER_6_194 VSS VDD scs8hd_fill_1
XFILLER_8_66 VSS VDD scs8hd_decap_4
XFILLER_40_3 VDD VSS scs8hd_fill_2
XANTENNA__673__D _572_/X VSS VDD scs8hd_diode_2
X_580_ _580_/A _578_/X _580_/X VSS VDD scs8hd_xor2_4
XPHY_255 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_244 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_233 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_222 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_52 VDD VSS scs8hd_fill_2
XPHY_211 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_200 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_17_75 VDD VSS scs8hd_fill_2
XFILLER_33_96 VDD VSS scs8hd_fill_2
XANTENNA__401__A _401_/A VSS VDD scs8hd_diode_2
XFILLER_30_252 VSS VDD scs8hd_fill_1
XFILLER_22_219 VSS VDD scs8hd_fill_1
XANTENNA__668__D _551_/X VSS VDD scs8hd_diode_2
XANTENNA__696__RESETB _350_/X VSS VDD scs8hd_diode_2
XFILLER_21_230 VDD VSS scs8hd_fill_2
XFILLER_0_156 VSS VDD scs8hd_decap_12
XFILLER_0_101 VDD VSS scs8hd_fill_2
XFILLER_0_112 VSS VDD scs8hd_decap_4
XFILLER_0_134 VDD VSS scs8hd_fill_2
XFILLER_28_41 VSS VDD scs8hd_decap_4
XFILLER_28_30 VSS VDD scs8hd_fill_1
X_632_ _694_/Q _632_/Y VSS VDD scs8hd_inv_8
X_563_ _563_/A _566_/A VSS VDD scs8hd_buf_1
X_494_ _491_/X _492_/X _494_/X VSS VDD scs8hd_xor2_4
XFILLER_8_212 VDD VSS scs8hd_fill_2
XFILLER_8_245 VSS VDD scs8hd_decap_8
XFILLER_12_252 VSS VDD scs8hd_fill_1
XANTENNA__543__A2N _539_/Y VSS VDD scs8hd_diode_2
XFILLER_5_67 VDD VSS scs8hd_fill_2
XFILLER_5_34 VDD VSS scs8hd_fill_2
XFILLER_39_116 VDD VSS scs8hd_fill_2
XFILLER_14_32 VDD VSS scs8hd_fill_2
XFILLER_14_43 VDD VSS scs8hd_fill_2
XFILLER_5_215 VSS VDD scs8hd_fill_1
XFILLER_5_237 VSS VDD scs8hd_decap_6
XFILLER_39_95 VDD VSS scs8hd_fill_2
XFILLER_39_62 VDD VSS scs8hd_fill_2
X_546_ _546_/A _546_/Y VSS VDD scs8hd_inv_8
XFILLER_29_193 VDD VSS scs8hd_fill_2
X_615_ _610_/Y _611_/Y _616_/A _616_/B _685_/D VSS VDD scs8hd_a2bb2o_4
X_477_ _476_/X _477_/X VSS VDD scs8hd_buf_1
XANTENNA__644__RESETB _413_/X VSS VDD scs8hd_diode_2
XFILLER_35_174 VSS VDD scs8hd_fill_1
XFILLER_35_152 VSS VDD scs8hd_decap_8
XANTENNA__681__D _600_/X VSS VDD scs8hd_diode_2
XPHY_64 VSS VDD scs8hd_decap_3
XPHY_53 VSS VDD scs8hd_decap_3
XFILLER_25_53 VDD VSS scs8hd_fill_2
X_331_ _605_/A x[28] _331_/X VSS VDD scs8hd_and2_4
X_400_ _401_/A _400_/X VSS VDD scs8hd_buf_1
XPHY_20 VSS VDD scs8hd_decap_3
XPHY_31 VSS VDD scs8hd_decap_3
XPHY_42 VSS VDD scs8hd_decap_3
XFILLER_41_177 VDD VSS scs8hd_fill_2
XPHY_75 VSS VDD scs8hd_decap_3
XPHY_97 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_86 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_37_9 VDD VSS scs8hd_fill_2
XFILLER_1_240 VSS VDD scs8hd_decap_4
X_529_ _524_/Y _525_/Y _527_/X _528_/X _661_/D VSS VDD scs8hd_a2bb2o_4
XANTENNA__348__B2 _347_/X VSS VDD scs8hd_diode_2
XFILLER_17_174 VSS VDD scs8hd_decap_4
XANTENNA__676__D _580_/X VSS VDD scs8hd_diode_2
XANTENNA__578__A1 _574_/Y VSS VDD scs8hd_diode_2
XANTENNA__578__B2 _678_/Q VSS VDD scs8hd_diode_2
XANTENNA__404__A _405_/A VSS VDD scs8hd_diode_2
XANTENNA__634__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_37_236 VDD VSS scs8hd_fill_2
XFILLER_20_125 VDD VSS scs8hd_fill_2
XFILLER_9_181 VDD VSS scs8hd_fill_2
XFILLER_28_203 VSS VDD scs8hd_decap_6
XFILLER_22_54 VSS VDD scs8hd_fill_1
XANTENNA__657__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_22_43 VSS VDD scs8hd_decap_4
XFILLER_22_32 VDD VSS scs8hd_fill_2
XFILLER_7_118 VSS VDD scs8hd_decap_4
XFILLER_0_3 VSS VDD scs8hd_decap_6
XFILLER_19_214 VDD VSS scs8hd_fill_2
XFILLER_19_225 VDD VSS scs8hd_fill_2
XFILLER_19_236 VSS VDD scs8hd_decap_8
XFILLER_6_162 VSS VDD scs8hd_decap_6
XFILLER_33_3 VSS VDD scs8hd_decap_4
XFILLER_25_217 VDD VSS scs8hd_fill_2
XANTENNA__692__RESETB _355_/X VSS VDD scs8hd_diode_2
XANTENNA__478__B1 _473_/A VSS VDD scs8hd_diode_2
XPHY_256 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_245 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_234 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_223 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_42 VSS VDD scs8hd_decap_4
XFILLER_31_209 VSS VDD scs8hd_decap_6
XPHY_212 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_201 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_24_250 VSS VDD scs8hd_decap_3
XFILLER_3_154 VDD VSS scs8hd_fill_2
XFILLER_3_110 VDD VSS scs8hd_fill_2
XFILLER_3_176 VSS VDD scs8hd_decap_3
XANTENNA__639__RESETB _419_/X VSS VDD scs8hd_diode_2
XANTENNA__684__D _684_/D VSS VDD scs8hd_diode_2
XFILLER_0_168 VSS VDD scs8hd_decap_12
XFILLER_0_146 VDD VSS scs8hd_fill_2
XANTENNA__502__A _502_/A VSS VDD scs8hd_diode_2
X_493_ _488_/Y _489_/Y _491_/X _492_/X _493_/X VSS VDD scs8hd_a2bb2o_4
X_631_ _691_/Q _631_/Y VSS VDD scs8hd_inv_8
X_562_ _597_/A x[18] _563_/A VSS VDD scs8hd_and2_4
XFILLER_8_202 VSS VDD scs8hd_fill_1
XANTENNA__543__A1N _538_/Y VSS VDD scs8hd_diode_2
XANTENNA__412__A _410_/A VSS VDD scs8hd_diode_2
XANTENNA__640__RESETB _418_/X VSS VDD scs8hd_diode_2
XANTENNA__614__B1 _685_/Q VSS VDD scs8hd_diode_2
XANTENNA__679__D _593_/X VSS VDD scs8hd_diode_2
XFILLER_38_194 VDD VSS scs8hd_fill_2
XFILLER_30_98 VDD VSS scs8hd_fill_2
XFILLER_30_32 VSS VDD scs8hd_decap_3
XFILLER_39_41 VDD VSS scs8hd_fill_2
XFILLER_29_172 VSS VDD scs8hd_decap_8
X_545_ _545_/A _545_/Y VSS VDD scs8hd_inv_8
X_476_ _476_/A x[6] _476_/X VSS VDD scs8hd_and2_4
XANTENNA__407__A _405_/A VSS VDD scs8hd_diode_2
X_614_ _610_/Y _611_/Y _685_/Q _611_/A _616_/B VSS VDD scs8hd_o22a_4
XFILLER_35_120 VDD VSS scs8hd_fill_2
XANTENNA__690__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_41_123 VDD VSS scs8hd_fill_2
XFILLER_41_101 VSS VDD scs8hd_decap_4
XPHY_76 VSS VDD scs8hd_decap_3
XPHY_65 VSS VDD scs8hd_decap_3
XPHY_54 VSS VDD scs8hd_decap_3
XPHY_43 VSS VDD scs8hd_decap_3
XPHY_10 VSS VDD scs8hd_decap_3
XPHY_98 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_87 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_21 VSS VDD scs8hd_decap_3
XPHY_32 VSS VDD scs8hd_decap_3
XFILLER_41_97 VDD VSS scs8hd_fill_2
XFILLER_41_86 VSS VDD scs8hd_decap_4
XFILLER_41_53 VDD VSS scs8hd_fill_2
XFILLER_41_42 VDD VSS scs8hd_fill_2
XFILLER_41_31 VDD VSS scs8hd_fill_2
XFILLER_2_36 VSS VDD scs8hd_fill_1
XFILLER_32_189 VSS VDD scs8hd_decap_4
X_528_ _524_/Y _525_/Y _661_/Q _664_/Q _528_/X VSS VDD scs8hd_o22a_4
X_459_ _643_/Q _459_/Y VSS VDD scs8hd_inv_8
XFILLER_23_123 VDD VSS scs8hd_fill_2
XFILLER_23_101 VSS VDD scs8hd_decap_12
XANTENNA__692__D _692_/D VSS VDD scs8hd_diode_2
XFILLER_11_12 VDD VSS scs8hd_fill_2
XFILLER_11_23 VDD VSS scs8hd_fill_2
XFILLER_11_56 VSS VDD scs8hd_fill_1
XANTENNA__510__A _660_/Q VSS VDD scs8hd_diode_2
XANTENNA__687__RESETB _362_/X VSS VDD scs8hd_diode_2
XANTENNA__578__A2 _575_/Y VSS VDD scs8hd_diode_2
XFILLER_36_75 VSS VDD scs8hd_decap_6
XFILLER_14_167 VSS VDD scs8hd_fill_1
XFILLER_37_215 VSS VDD scs8hd_fill_1
XFILLER_35_7 VDD VSS scs8hd_fill_2
XANTENNA__420__A _417_/A VSS VDD scs8hd_diode_2
XANTENNA__579__A2N _575_/Y VSS VDD scs8hd_diode_2
XFILLER_20_148 VSS VDD scs8hd_fill_1
XFILLER_28_215 VDD VSS scs8hd_fill_2
XANTENNA__687__D _687_/D VSS VDD scs8hd_diode_2
XFILLER_22_77 VSS VDD scs8hd_decap_3
XANTENNA__505__A _504_/X VSS VDD scs8hd_diode_2
XFILLER_34_207 VSS VDD scs8hd_decap_3
XFILLER_8_79 VSS VDD scs8hd_decap_12
XANTENNA__415__A _410_/A VSS VDD scs8hd_diode_2
XFILLER_6_174 VDD VSS scs8hd_fill_2
XFILLER_26_3 VDD VSS scs8hd_fill_2
XANTENNA__635__RESETB _423_/X VSS VDD scs8hd_diode_2
XANTENNA__478__B2 _474_/A VSS VDD scs8hd_diode_2
XANTENNA__478__A1 _473_/Y VSS VDD scs8hd_diode_2
XFILLER_17_66 VSS VDD scs8hd_decap_6
XFILLER_17_99 VDD VSS scs8hd_fill_2
XPHY_257 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_246 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_235 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_224 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_213 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_202 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_15_240 VSS VDD scs8hd_decap_4
XANTENNA__647__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_0_91 VDD VSS scs8hd_fill_2
XFILLER_28_32 VDD VSS scs8hd_fill_2
XFILLER_0_125 VDD VSS scs8hd_fill_2
X_630_ _627_/X _630_/B _630_/X VSS VDD scs8hd_xor2_4
X_492_ _488_/Y _489_/Y _488_/A _489_/A _492_/X VSS VDD scs8hd_o22a_4
XFILLER_28_98 VDD VSS scs8hd_fill_2
XFILLER_28_87 VSS VDD scs8hd_fill_1
XFILLER_28_76 VSS VDD scs8hd_decap_4
X_561_ _518_/A _597_/A VSS VDD scs8hd_buf_1
XFILLER_39_107 VSS VDD scs8hd_decap_3
XFILLER_5_47 VDD VSS scs8hd_fill_2
XANTENNA__614__A1 _610_/Y VSS VDD scs8hd_diode_2
XANTENNA__614__B2 _611_/A VSS VDD scs8hd_diode_2
XANTENNA__550__B1 _548_/X VSS VDD scs8hd_diode_2
XANTENNA__603__A _603_/A VSS VDD scs8hd_diode_2
XFILLER_38_184 VSS VDD scs8hd_decap_4
XFILLER_38_151 VDD VSS scs8hd_fill_2
XFILLER_38_140 VDD VSS scs8hd_fill_2
XANTENNA__695__D _348_/X VSS VDD scs8hd_diode_2
XFILLER_30_11 VSS VDD scs8hd_decap_3
XFILLER_14_23 VDD VSS scs8hd_fill_2
XFILLER_30_66 VSS VDD scs8hd_decap_4
XFILLER_39_86 VSS VDD scs8hd_decap_6
XFILLER_29_184 VDD VSS scs8hd_fill_2
X_613_ _612_/X _616_/A VSS VDD scs8hd_buf_1
X_544_ _544_/A _544_/B _544_/X VSS VDD scs8hd_xor2_4
X_475_ _518_/A _476_/A VSS VDD scs8hd_buf_1
XANTENNA__423__A _366_/A VSS VDD scs8hd_diode_2
XANTENNA__599__B1 _595_/A VSS VDD scs8hd_diode_2
XFILLER_35_165 VSS VDD scs8hd_decap_3
XPHY_77 VSS VDD scs8hd_decap_3
XPHY_66 VSS VDD scs8hd_decap_3
XPHY_55 VSS VDD scs8hd_decap_3
XFILLER_26_198 VSS VDD scs8hd_decap_8
XFILLER_26_154 VDD VSS scs8hd_fill_2
XFILLER_26_132 VDD VSS scs8hd_fill_2
XANTENNA__508__A _508_/A VSS VDD scs8hd_diode_2
XFILLER_25_33 VDD VSS scs8hd_fill_2
XPHY_44 VSS VDD scs8hd_decap_3
XPHY_99 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_88 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_11 VSS VDD scs8hd_decap_3
XPHY_22 VSS VDD scs8hd_decap_3
XPHY_33 VSS VDD scs8hd_decap_3
XANTENNA__683__RESETB _367_/X VSS VDD scs8hd_diode_2
XANTENNA__514__B1 _515_/A VSS VDD scs8hd_diode_2
XFILLER_2_26 VSS VDD scs8hd_fill_1
XFILLER_2_15 VSS VDD scs8hd_decap_4
X_527_ _527_/A _527_/X VSS VDD scs8hd_buf_1
XANTENNA__418__A _417_/A VSS VDD scs8hd_diode_2
XFILLER_17_132 VSS VDD scs8hd_decap_4
XFILLER_17_143 VDD VSS scs8hd_fill_2
X_389_ _389_/A _389_/X VSS VDD scs8hd_buf_1
XFILLER_32_146 VSS VDD scs8hd_decap_6
X_458_ _458_/A _456_/X _458_/X VSS VDD scs8hd_xor2_4
XFILLER_23_113 VSS VDD scs8hd_fill_1
XFILLER_36_87 VSS VDD scs8hd_fill_1
XFILLER_36_32 VDD VSS scs8hd_fill_2
XANTENNA__500__A2N _496_/Y VSS VDD scs8hd_diode_2
XFILLER_14_102 VSS VDD scs8hd_decap_12
XFILLER_14_135 VDD VSS scs8hd_fill_2
XFILLER_28_7 VSS VDD scs8hd_decap_4
XANTENNA__579__A1N _574_/Y VSS VDD scs8hd_diode_2
XANTENNA__680__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__611__A _611_/A VSS VDD scs8hd_diode_2
XFILLER_22_23 VDD VSS scs8hd_fill_2
XFILLER_7_109 VDD VSS scs8hd_fill_2
XFILLER_11_138 VSS VDD scs8hd_fill_1
XFILLER_42_230 VSS VDD scs8hd_fill_1
XFILLER_8_25 VDD VSS scs8hd_fill_2
XFILLER_10_193 VSS VDD scs8hd_decap_4
XANTENNA__431__A _431_/A VSS VDD scs8hd_diode_2
XFILLER_6_186 VDD VSS scs8hd_fill_2
XFILLER_19_3 VDD VSS scs8hd_fill_2
XANTENNA__606__A _605_/X VSS VDD scs8hd_diode_2
XANTENNA__478__A2 _474_/Y VSS VDD scs8hd_diode_2
XPHY_225 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_214 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_203 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_16_208 VDD VSS scs8hd_fill_2
XPHY_258 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_247 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_236 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__516__A _516_/A VSS VDD scs8hd_diode_2
XFILLER_3_123 VDD VSS scs8hd_fill_2
XFILLER_3_101 VDD VSS scs8hd_fill_2
XANTENNA__426__A _633_/Q VSS VDD scs8hd_diode_2
XANTENNA__336__A _693_/Q VSS VDD scs8hd_diode_2
XFILLER_28_22 VDD VSS scs8hd_fill_2
XFILLER_28_11 VSS VDD scs8hd_fill_1
X_560_ _560_/A _560_/Y VSS VDD scs8hd_inv_8
X_491_ _490_/X _491_/X VSS VDD scs8hd_buf_1
XFILLER_12_244 VSS VDD scs8hd_decap_8
XFILLER_8_215 VSS VDD scs8hd_decap_3
XFILLER_5_59 VDD VSS scs8hd_fill_2
XANTENNA__678__RESETB _372_/X VSS VDD scs8hd_diode_2
XFILLER_10_7 VDD VSS scs8hd_fill_2
X_689_ _681_/CLK _629_/X _624_/A _360_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__614__A2 _611_/Y VSS VDD scs8hd_diode_2
XANTENNA__550__B2 _551_/B VSS VDD scs8hd_diode_2
XFILLER_30_45 VSS VDD scs8hd_fill_1
XFILLER_30_23 VSS VDD scs8hd_decap_8
XFILLER_5_218 VDD VSS scs8hd_fill_2
X_543_ _538_/Y _539_/Y _544_/A _544_/B _543_/X VSS VDD scs8hd_a2bb2o_4
X_612_ _605_/A x[25] _612_/X VSS VDD scs8hd_and2_4
X_474_ _474_/A _474_/Y VSS VDD scs8hd_inv_8
XANTENNA__637__CLK _648_/CLK VSS VDD scs8hd_diode_2
XANTENNA__599__A1 _595_/Y VSS VDD scs8hd_diode_2
XANTENNA__599__B2 _684_/Q VSS VDD scs8hd_diode_2
XFILLER_35_177 VDD VSS scs8hd_fill_2
XFILLER_6_91 VSS VDD scs8hd_fill_1
XFILLER_26_144 VSS VDD scs8hd_decap_4
XPHY_12 VSS VDD scs8hd_decap_3
XFILLER_41_136 VSS VDD scs8hd_decap_3
XFILLER_41_114 VSS VDD scs8hd_decap_4
XPHY_78 VSS VDD scs8hd_decap_3
XPHY_67 VSS VDD scs8hd_decap_3
XPHY_56 VSS VDD scs8hd_decap_3
XFILLER_26_188 VDD VSS scs8hd_fill_2
XANTENNA__508__B _508_/B VSS VDD scs8hd_diode_2
XFILLER_25_89 VSS VDD scs8hd_decap_4
XPHY_45 VSS VDD scs8hd_decap_3
XPHY_89 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_23 VSS VDD scs8hd_decap_3
XPHY_34 VSS VDD scs8hd_decap_3
XFILLER_41_66 VSS VDD scs8hd_fill_1
XANTENNA__524__A _661_/Q VSS VDD scs8hd_diode_2
XANTENNA__514__B2 _513_/X VSS VDD scs8hd_diode_2
XFILLER_1_232 VDD VSS scs8hd_fill_2
X_526_ _547_/A x[13] _527_/A VSS VDD scs8hd_and2_4
XANTENNA__450__B1 _451_/A VSS VDD scs8hd_diode_2
X_388_ _402_/A _389_/A VSS VDD scs8hd_buf_1
XANTENNA__434__A _434_/A VSS VDD scs8hd_diode_2
X_457_ _452_/Y _453_/Y _458_/A _456_/X _457_/X VSS VDD scs8hd_a2bb2o_4
XANTENNA__609__A _609_/A VSS VDD scs8hd_diode_2
XFILLER_23_158 VDD VSS scs8hd_fill_2
XANTENNA__344__A _344_/A VSS VDD scs8hd_diode_2
XFILLER_36_11 VSS VDD scs8hd_decap_3
XANTENNA__500__A1N _495_/Y VSS VDD scs8hd_diode_2
XANTENNA__432__B1 _633_/Q VSS VDD scs8hd_diode_2
XFILLER_14_114 VSS VDD scs8hd_decap_4
XFILLER_14_125 VSS VDD scs8hd_decap_3
XANTENNA__519__A _547_/A VSS VDD scs8hd_diode_2
XFILLER_14_147 VDD VSS scs8hd_fill_2
XANTENNA__499__B1 _653_/Q VSS VDD scs8hd_diode_2
XANTENNA__429__A _518_/A VSS VDD scs8hd_diode_2
X_509_ _657_/Q _509_/Y VSS VDD scs8hd_inv_8
XFILLER_9_184 VDD VSS scs8hd_fill_2
XANTENNA__339__A _339_/A VSS VDD scs8hd_diode_2
XFILLER_22_57 VDD VSS scs8hd_fill_2
XFILLER_11_117 VSS VDD scs8hd_fill_1
XFILLER_11_128 VDD VSS scs8hd_fill_2
XANTENNA__348__A2N _344_/Y VSS VDD scs8hd_diode_2
XFILLER_6_154 VDD VSS scs8hd_fill_2
XFILLER_12_90 VDD VSS scs8hd_fill_2
XFILLER_6_198 VSS VDD scs8hd_decap_4
XFILLER_25_209 VDD VSS scs8hd_fill_2
XPHY_259 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_248 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_237 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_226 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_34 VDD VSS scs8hd_fill_2
XPHY_215 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_204 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_24_242 VSS VDD scs8hd_decap_8
XFILLER_17_79 VDD VSS scs8hd_fill_2
XANTENNA__532__A _666_/Q VSS VDD scs8hd_diode_2
XFILLER_33_67 VDD VSS scs8hd_fill_2
XFILLER_33_56 VSS VDD scs8hd_decap_4
XANTENNA__670__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_30_212 VDD VSS scs8hd_fill_2
XANTENNA__437__B1N _436_/X VSS VDD scs8hd_diode_2
XANTENNA__674__RESETB _378_/X VSS VDD scs8hd_diode_2
XFILLER_31_3 VDD VSS scs8hd_fill_2
XANTENNA__617__A _687_/Q VSS VDD scs8hd_diode_2
XFILLER_0_71 VSS VDD scs8hd_decap_12
XFILLER_21_245 VSS VDD scs8hd_decap_8
XFILLER_21_234 VDD VSS scs8hd_fill_2
XANTENNA__693__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__352__A _373_/A VSS VDD scs8hd_diode_2
XFILLER_0_105 VSS VDD scs8hd_decap_4
XFILLER_0_138 VDD VSS scs8hd_fill_2
XANTENNA__CTS_buf_1_32_A _CTS_root/X VSS VDD scs8hd_diode_2
XANTENNA__608__B1 _609_/A VSS VDD scs8hd_diode_2
XFILLER_28_45 VSS VDD scs8hd_fill_1
X_490_ _476_/A x[8] _490_/X VSS VDD scs8hd_and2_4
XANTENNA__536__A2N _532_/Y VSS VDD scs8hd_diode_2
XANTENNA__527__A _527_/A VSS VDD scs8hd_diode_2
XFILLER_5_38 VDD VSS scs8hd_fill_2
XFILLER_5_27 VSS VDD scs8hd_decap_4
X_688_ _681_/CLK _688_/D _611_/A _361_/X VSS VDD scs8hd_dfrtp_4
XFILLER_14_47 VDD VSS scs8hd_fill_2
XFILLER_39_99 VDD VSS scs8hd_fill_2
XFILLER_39_55 VDD VSS scs8hd_fill_2
XFILLER_39_11 VSS VDD scs8hd_decap_4
X_542_ _538_/Y _539_/Y _538_/A _539_/A _544_/B VSS VDD scs8hd_o22a_4
XFILLER_29_197 VSS VDD scs8hd_decap_3
X_473_ _473_/A _473_/Y VSS VDD scs8hd_inv_8
X_611_ _611_/A _611_/Y VSS VDD scs8hd_inv_8
XFILLER_20_90 VDD VSS scs8hd_fill_2
XANTENNA__599__A2 _596_/Y VSS VDD scs8hd_diode_2
XFILLER_35_123 VDD VSS scs8hd_fill_2
XANTENNA__630__A _627_/X VSS VDD scs8hd_diode_2
XPHY_46 VSS VDD scs8hd_decap_3
XPHY_13 VSS VDD scs8hd_decap_3
XPHY_24 VSS VDD scs8hd_decap_3
XPHY_35 VSS VDD scs8hd_decap_3
XPHY_79 VSS VDD scs8hd_decap_3
XPHY_68 VSS VDD scs8hd_decap_3
XPHY_57 VSS VDD scs8hd_decap_3
XFILLER_25_57 VSS VDD scs8hd_decap_4
XANTENNA__540__A _547_/A VSS VDD scs8hd_diode_2
XFILLER_1_200 VDD VSS scs8hd_fill_2
XFILLER_9_3 VDD VSS scs8hd_fill_2
XFILLER_32_104 VSS VDD scs8hd_decap_6
X_525_ _664_/Q _525_/Y VSS VDD scs8hd_inv_8
XANTENNA__450__B2 _449_/X VSS VDD scs8hd_diode_2
X_456_ _452_/Y _453_/Y _452_/A _644_/Q _456_/X VSS VDD scs8hd_o22a_4
XFILLER_17_123 VDD VSS scs8hd_fill_2
XFILLER_17_178 VSS VDD scs8hd_fill_1
XFILLER_40_181 VSS VDD scs8hd_fill_1
X_387_ _386_/A _387_/X VSS VDD scs8hd_buf_1
XANTENNA__434__B _434_/B VSS VDD scs8hd_diode_2
XANTENNA__609__B _609_/B VSS VDD scs8hd_diode_2
XFILLER_31_181 VDD VSS scs8hd_fill_2
XANTENNA__625__A _625_/A VSS VDD scs8hd_diode_2
XANTENNA__360__A _363_/A VSS VDD scs8hd_diode_2
XFILLER_11_59 VDD VSS scs8hd_fill_2
XFILLER_36_23 VDD VSS scs8hd_fill_2
XANTENNA__432__B2 _638_/Q VSS VDD scs8hd_diode_2
XANTENNA__432__A1 _426_/Y VSS VDD scs8hd_diode_2
XANTENNA__519__B x[12] VSS VDD scs8hd_diode_2
XANTENNA__499__B2 _496_/A VSS VDD scs8hd_diode_2
XANTENNA__499__A1 _495_/Y VSS VDD scs8hd_diode_2
XFILLER_37_218 VDD VSS scs8hd_fill_2
X_508_ _508_/A _508_/B _508_/X VSS VDD scs8hd_xor2_4
X_439_ _640_/Q _439_/Y VSS VDD scs8hd_inv_8
XANTENNA__445__A _445_/A VSS VDD scs8hd_diode_2
XFILLER_13_192 VDD VSS scs8hd_fill_2
XFILLER_20_118 VSS VDD scs8hd_decap_4
XFILLER_20_129 VDD VSS scs8hd_fill_2
XFILLER_9_163 VDD VSS scs8hd_fill_2
XFILLER_9_174 VSS VDD scs8hd_decap_4
XANTENNA__669__RESETB _384_/X VSS VDD scs8hd_diode_2
XFILLER_36_251 VDD VSS scs8hd_fill_2
XFILLER_22_47 VSS VDD scs8hd_fill_1
XANTENNA__355__A _357_/A VSS VDD scs8hd_diode_2
XANTENNA__348__A1N _343_/Y VSS VDD scs8hd_diode_2
XFILLER_8_38 VDD VSS scs8hd_fill_2
XANTENNA__341__B1 _339_/X VSS VDD scs8hd_diode_2
XFILLER_6_144 VSS VDD scs8hd_decap_4
XFILLER_10_151 VDD VSS scs8hd_fill_2
XFILLER_12_80 VSS VDD scs8hd_fill_1
XANTENNA__670__RESETB _383_/X VSS VDD scs8hd_diode_2
XFILLER_33_232 VSS VDD scs8hd_decap_12
XFILLER_18_251 VDD VSS scs8hd_fill_2
XFILLER_17_25 VDD VSS scs8hd_fill_2
XPHY_249 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_238 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_227 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_216 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_205 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_24_210 VSS VDD scs8hd_decap_4
XFILLER_17_58 VSS VDD scs8hd_decap_3
XFILLER_3_114 VDD VSS scs8hd_fill_2
XANTENNA__571__B1 _673_/Q VSS VDD scs8hd_diode_2
XFILLER_15_221 VSS VDD scs8hd_decap_4
XFILLER_15_232 VDD VSS scs8hd_fill_2
XFILLER_30_202 VDD VSS scs8hd_fill_2
XFILLER_24_3 VDD VSS scs8hd_fill_2
XFILLER_0_61 VSS VDD scs8hd_fill_1
XFILLER_0_83 VSS VDD scs8hd_decap_8
XFILLER_0_94 VSS VDD scs8hd_decap_4
XANTENNA__608__B2 _609_/B VSS VDD scs8hd_diode_2
XANTENNA__536__A1N _531_/Y VSS VDD scs8hd_diode_2
XFILLER_8_206 VSS VDD scs8hd_decap_4
XFILLER_12_202 VSS VDD scs8hd_decap_12
X_687_ _681_/CLK _687_/D _687_/Q _362_/X VSS VDD scs8hd_dfrtp_4
XFILLER_18_90 VDD VSS scs8hd_fill_2
XANTENNA__535__B1 _663_/Q VSS VDD scs8hd_diode_2
XANTENNA__453__A _644_/Q VSS VDD scs8hd_diode_2
XFILLER_38_198 VDD VSS scs8hd_fill_2
XFILLER_38_154 VDD VSS scs8hd_fill_2
XFILLER_38_132 VDD VSS scs8hd_fill_2
XFILLER_38_110 VSS VDD scs8hd_decap_4
XANTENNA__363__A _363_/A VSS VDD scs8hd_diode_2
XANTENNA__660__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_5_209 VSS VDD scs8hd_decap_6
XFILLER_39_78 VDD VSS scs8hd_fill_2
XFILLER_39_45 VDD VSS scs8hd_fill_2
XFILLER_29_143 VDD VSS scs8hd_fill_2
XFILLER_29_121 VSS VDD scs8hd_fill_1
X_610_ _685_/Q _610_/Y VSS VDD scs8hd_inv_8
XANTENNA__538__A _538_/A VSS VDD scs8hd_diode_2
X_541_ _540_/X _544_/A VSS VDD scs8hd_buf_1
X_472_ _469_/X _470_/X _472_/X VSS VDD scs8hd_xor2_4
XFILLER_35_113 VSS VDD scs8hd_decap_4
XANTENNA__683__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__448__A _448_/A VSS VDD scs8hd_diode_2
XFILLER_6_93 VSS VDD scs8hd_decap_3
XANTENNA__630__B _630_/B VSS VDD scs8hd_diode_2
XPHY_69 VSS VDD scs8hd_decap_3
XPHY_58 VSS VDD scs8hd_decap_3
XFILLER_26_179 VSS VDD scs8hd_decap_3
XPHY_47 VSS VDD scs8hd_decap_3
XANTENNA__358__A _373_/A VSS VDD scs8hd_diode_2
XPHY_14 VSS VDD scs8hd_decap_3
XPHY_25 VSS VDD scs8hd_decap_3
XPHY_36 VSS VDD scs8hd_decap_3
XFILLER_41_57 VSS VDD scs8hd_decap_4
XANTENNA__540__B x[15] VSS VDD scs8hd_diode_2
XFILLER_1_245 VSS VDD scs8hd_decap_8
XFILLER_2_29 VDD VSS scs8hd_fill_2
X_386_ _386_/A _386_/X VSS VDD scs8hd_buf_1
X_524_ _661_/Q _524_/Y VSS VDD scs8hd_inv_8
XFILLER_15_91 VDD VSS scs8hd_fill_2
X_455_ _454_/X _458_/A VSS VDD scs8hd_buf_1
XFILLER_23_116 VDD VSS scs8hd_fill_2
XANTENNA__665__RESETB _389_/X VSS VDD scs8hd_diode_2
XFILLER_31_171 VDD VSS scs8hd_fill_2
XFILLER_31_160 VDD VSS scs8hd_fill_2
XFILLER_11_16 VSS VDD scs8hd_decap_4
XFILLER_11_27 VDD VSS scs8hd_fill_2
XANTENNA__432__A2 _427_/Y VSS VDD scs8hd_diode_2
XANTENNA__551__A _548_/X VSS VDD scs8hd_diode_2
XANTENNA__499__A2 _496_/Y VSS VDD scs8hd_diode_2
X_CTS_buf_1_32 _CTS_root/X _667_/CLK VSS VDD scs8hd_clkbuf_4
X_369_ _370_/A _369_/X VSS VDD scs8hd_buf_1
XFILLER_26_90 VDD VSS scs8hd_fill_2
X_507_ _502_/Y _503_/Y _508_/A _508_/B _507_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_9_120 VDD VSS scs8hd_fill_2
XFILLER_9_131 VDD VSS scs8hd_fill_2
X_438_ _438_/A _438_/Y VSS VDD scs8hd_inv_8
XFILLER_13_182 VSS VDD scs8hd_fill_1
XANTENNA__461__A _461_/A VSS VDD scs8hd_diode_2
XFILLER_28_219 VDD VSS scs8hd_fill_2
XANTENNA__371__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_42_211 VSS VDD scs8hd_decap_6
XFILLER_19_219 VSS VDD scs8hd_decap_4
XANTENNA__546__A _546_/A VSS VDD scs8hd_diode_2
XANTENNA__341__B2 _340_/X VSS VDD scs8hd_diode_2
XFILLER_6_178 VDD VSS scs8hd_fill_2
XFILLER_26_7 VSS VDD scs8hd_decap_4
XPHY_239 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_228 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_217 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_206 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__366__A _366_/A VSS VDD scs8hd_diode_2
XFILLER_3_148 VSS VDD scs8hd_decap_4
XANTENNA__571__A1 _567_/Y VSS VDD scs8hd_diode_2
XANTENNA__571__B2 _676_/Q VSS VDD scs8hd_diode_2
XFILLER_23_91 VSS VDD scs8hd_decap_8
XFILLER_17_3 VDD VSS scs8hd_fill_2
XFILLER_9_71 VDD VSS scs8hd_fill_2
XFILLER_28_14 VDD VSS scs8hd_fill_2
XFILLER_0_118 VDD VSS scs8hd_fill_2
XFILLER_34_90 VDD VSS scs8hd_fill_2
X_686_ _681_/CLK _686_/D _603_/A _363_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__535__B2 _666_/Q VSS VDD scs8hd_diode_2
XANTENNA__535__A1 _531_/Y VSS VDD scs8hd_diode_2
XFILLER_7_240 VSS VDD scs8hd_decap_4
XFILLER_38_144 VSS VDD scs8hd_decap_4
XANTENNA__471__B1 _469_/X VSS VDD scs8hd_diode_2
XFILLER_14_27 VSS VDD scs8hd_decap_4
XFILLER_30_37 VDD VSS scs8hd_fill_2
X_540_ _547_/A x[15] _540_/X VSS VDD scs8hd_and2_4
XFILLER_29_111 VDD VSS scs8hd_fill_2
XANTENNA__554__A _547_/A VSS VDD scs8hd_diode_2
X_471_ _466_/Y _467_/Y _469_/X _470_/X _471_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_4_221 VDD VSS scs8hd_fill_2
XFILLER_20_81 VSS VDD scs8hd_decap_6
X_669_ _667_/CLK _669_/D _552_/A _384_/X VSS VDD scs8hd_dfrtp_4
XFILLER_6_61 VDD VSS scs8hd_fill_2
XFILLER_6_83 VSS VDD scs8hd_decap_8
XANTENNA__661__RESETB _393_/X VSS VDD scs8hd_diode_2
XPHY_59 VSS VDD scs8hd_decap_3
XFILLER_26_136 VDD VSS scs8hd_fill_2
XANTENNA__374__A _402_/A VSS VDD scs8hd_diode_2
XFILLER_25_37 VDD VSS scs8hd_fill_2
XPHY_48 VSS VDD scs8hd_decap_3
XPHY_15 VSS VDD scs8hd_decap_3
XPHY_26 VSS VDD scs8hd_decap_3
XPHY_37 VSS VDD scs8hd_decap_3
XFILLER_41_69 VDD VSS scs8hd_fill_2
XFILLER_41_36 VSS VDD scs8hd_decap_4
XFILLER_2_19 VSS VDD scs8hd_fill_1
XFILLER_1_224 VDD VSS scs8hd_fill_2
XFILLER_17_103 VSS VDD scs8hd_decap_4
XFILLER_17_114 VDD VSS scs8hd_fill_2
XFILLER_17_147 VSS VDD scs8hd_decap_4
X_523_ _520_/X _521_/X _660_/D VSS VDD scs8hd_xor2_4
X_385_ _386_/A _385_/X VSS VDD scs8hd_buf_1
XFILLER_32_139 VSS VDD scs8hd_fill_1
X_454_ _461_/A x[3] _454_/X VSS VDD scs8hd_and2_4
XANTENNA__650__CLK _651_/CLK VSS VDD scs8hd_diode_2
XANTENNA__459__A _643_/Q VSS VDD scs8hd_diode_2
XFILLER_23_139 VDD VSS scs8hd_fill_2
XFILLER_36_36 VSS VDD scs8hd_decap_3
XANTENNA__369__A _370_/A VSS VDD scs8hd_diode_2
XFILLER_22_183 VSS VDD scs8hd_fill_1
XFILLER_14_139 VSS VDD scs8hd_decap_8
XANTENNA__551__B _551_/B VSS VDD scs8hd_diode_2
XANTENNA__673__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_26_80 VSS VDD scs8hd_fill_1
X_506_ _502_/Y _503_/Y _502_/A _658_/Q _508_/B VSS VDD scs8hd_o22a_4
X_368_ _370_/A _368_/X VSS VDD scs8hd_buf_1
X_437_ _635_/Q _435_/X _436_/X _437_/Y VSS VDD scs8hd_a21boi_4
XFILLER_13_161 VDD VSS scs8hd_fill_2
XFILLER_13_172 VSS VDD scs8hd_decap_4
XANTENNA__461__B x[4] VSS VDD scs8hd_diode_2
XFILLER_28_209 VSS VDD scs8hd_fill_1
XFILLER_3_95 VSS VDD scs8hd_decap_4
XFILLER_3_62 VSS VDD scs8hd_decap_4
XFILLER_11_109 VDD VSS scs8hd_fill_2
XFILLER_22_27 VSS VDD scs8hd_decap_4
XANTENNA__696__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_0_9 VSS VDD scs8hd_fill_1
XANTENNA__CTS_buf_1_48_A _CTS_root/X VSS VDD scs8hd_diode_2
XFILLER_19_209 VSS VDD scs8hd_decap_3
XFILLER_42_234 VDD VSS scs8hd_fill_2
XFILLER_27_231 VDD VSS scs8hd_fill_2
XFILLER_8_29 VDD VSS scs8hd_fill_2
XANTENNA__562__A _597_/A VSS VDD scs8hd_diode_2
XFILLER_33_9 VDD VSS scs8hd_fill_2
XANTENNA__629__B1 _627_/X VSS VDD scs8hd_diode_2
XFILLER_12_93 VDD VSS scs8hd_fill_2
XFILLER_33_245 VSS VDD scs8hd_decap_8
XANTENNA__472__A _469_/X VSS VDD scs8hd_diode_2
XPHY_207 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_229 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_48 VDD VSS scs8hd_fill_2
XPHY_218 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__382__A _386_/A VSS VDD scs8hd_diode_2
XANTENNA__571__A2 _568_/Y VSS VDD scs8hd_diode_2
XFILLER_30_215 VDD VSS scs8hd_fill_2
XFILLER_15_245 VDD VSS scs8hd_fill_2
XFILLER_2_171 VSS VDD scs8hd_fill_1
XFILLER_0_41 VDD VSS scs8hd_fill_2
XFILLER_0_63 VDD VSS scs8hd_fill_2
XANTENNA__467__A _648_/Q VSS VDD scs8hd_diode_2
XFILLER_21_215 VDD VSS scs8hd_fill_2
XFILLER_21_226 VDD VSS scs8hd_fill_2
XFILLER_28_48 VDD VSS scs8hd_fill_2
XFILLER_28_37 VDD VSS scs8hd_fill_2
XFILLER_28_26 VSS VDD scs8hd_decap_4
XFILLER_12_215 VSS VDD scs8hd_decap_6
XANTENNA__377__A _375_/A VSS VDD scs8hd_diode_2
XANTENNA__656__RESETB _399_/X VSS VDD scs8hd_diode_2
X_685_ _681_/CLK _685_/D _685_/Q _364_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__535__A2 _532_/Y VSS VDD scs8hd_diode_2
XANTENNA__471__B2 _470_/X VSS VDD scs8hd_diode_2
XFILLER_30_16 VSS VDD scs8hd_decap_4
XFILLER_29_189 VDD VSS scs8hd_fill_2
XFILLER_29_123 VSS VDD scs8hd_decap_12
XANTENNA__554__B x[17] VSS VDD scs8hd_diode_2
X_470_ _466_/Y _467_/Y _645_/Q _648_/Q _470_/X VSS VDD scs8hd_o22a_4
XFILLER_4_233 VSS VDD scs8hd_decap_3
XANTENNA__570__A _570_/A VSS VDD scs8hd_diode_2
XFILLER_29_80 VSS VDD scs8hd_decap_3
XFILLER_20_93 VDD VSS scs8hd_fill_2
X_668_ _667_/CLK _551_/X _539_/A _385_/X VSS VDD scs8hd_dfrtp_4
X_599_ _595_/Y _596_/Y _595_/A _684_/Q _601_/B VSS VDD scs8hd_o22a_4
XFILLER_35_148 VDD VSS scs8hd_fill_2
XANTENNA__480__A _477_/X VSS VDD scs8hd_diode_2
XFILLER_26_104 VSS VDD scs8hd_fill_1
XFILLER_34_192 VDD VSS scs8hd_fill_2
XFILLER_26_148 VSS VDD scs8hd_fill_1
XFILLER_25_27 VSS VDD scs8hd_decap_4
XPHY_49 VSS VDD scs8hd_decap_3
XPHY_16 VSS VDD scs8hd_decap_3
XANTENNA__572__A2N _568_/Y VSS VDD scs8hd_diode_2
XPHY_27 VSS VDD scs8hd_decap_3
XPHY_38 VSS VDD scs8hd_decap_3
XFILLER_41_15 VSS VDD scs8hd_decap_12
XANTENNA__390__A _389_/A VSS VDD scs8hd_diode_2
XFILLER_1_236 VDD VSS scs8hd_fill_2
X_453_ _644_/Q _453_/Y VSS VDD scs8hd_inv_8
X_522_ _516_/Y _517_/Y _520_/X _521_/X _522_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_40_184 VDD VSS scs8hd_fill_2
XFILLER_40_173 VDD VSS scs8hd_fill_2
XFILLER_40_151 VDD VSS scs8hd_fill_2
X_384_ _386_/A _384_/X VSS VDD scs8hd_buf_1
XFILLER_25_181 VDD VSS scs8hd_fill_2
XANTENNA__475__A _518_/A VSS VDD scs8hd_diode_2
XFILLER_31_184 VDD VSS scs8hd_fill_2
XANTENNA__385__A _386_/A VSS VDD scs8hd_diode_2
XFILLER_14_118 VSS VDD scs8hd_fill_1
XFILLER_22_151 VDD VSS scs8hd_fill_2
XFILLER_7_3 VSS VDD scs8hd_decap_3
X_436_ _635_/Q _435_/X _436_/X VSS VDD scs8hd_or2_4
X_505_ _504_/X _508_/A VSS VDD scs8hd_buf_1
XANTENNA__592__B1 _679_/Q VSS VDD scs8hd_diode_2
X_367_ _370_/A _367_/X VSS VDD scs8hd_buf_1
XFILLER_13_184 VDD VSS scs8hd_fill_2
XFILLER_3_52 VSS VDD scs8hd_decap_4
XFILLER_36_243 VSS VDD scs8hd_decap_8
XFILLER_42_246 VDD VSS scs8hd_fill_2
XFILLER_27_243 VSS VDD scs8hd_fill_1
XANTENNA__640__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_6_114 VDD VSS scs8hd_fill_2
XFILLER_6_158 VDD VSS scs8hd_fill_2
XFILLER_10_143 VSS VDD scs8hd_decap_6
XFILLER_10_154 VDD VSS scs8hd_fill_2
XFILLER_10_165 VDD VSS scs8hd_fill_2
XFILLER_12_50 VSS VDD scs8hd_fill_1
XFILLER_12_61 VDD VSS scs8hd_fill_2
XFILLER_12_72 VDD VSS scs8hd_fill_2
XANTENNA__562__B x[18] VSS VDD scs8hd_diode_2
XANTENNA__629__B2 _630_/B VSS VDD scs8hd_diode_2
XFILLER_37_91 VSS VDD scs8hd_decap_4
XFILLER_18_243 VSS VDD scs8hd_decap_8
XFILLER_33_224 VDD VSS scs8hd_fill_2
X_419_ _417_/A _419_/X VSS VDD scs8hd_buf_1
XANTENNA__472__B _470_/X VSS VDD scs8hd_diode_2
XANTENNA__565__B1 _566_/A VSS VDD scs8hd_diode_2
XANTENNA__663__CLK _651_/CLK VSS VDD scs8hd_diode_2
XPHY_219 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_208 VSS VDD scs8hd_tapvpwrvgnd_1
XFILLER_33_38 VDD VSS scs8hd_fill_2
XANTENNA__556__B1 _552_/A VSS VDD scs8hd_diode_2
XANTENNA__652__RESETB _404_/X VSS VDD scs8hd_diode_2
XFILLER_15_202 VDD VSS scs8hd_fill_2
XANTENNA__573__A _570_/X VSS VDD scs8hd_diode_2
XANTENNA__686__CLK _681_/CLK VSS VDD scs8hd_diode_2
XANTENNA__483__A _476_/A VSS VDD scs8hd_diode_2
XFILLER_21_238 VSS VDD scs8hd_decap_6
XANTENNA__633__D _633_/D VSS VDD scs8hd_diode_2
XFILLER_9_62 VSS VDD scs8hd_decap_3
XFILLER_9_95 VDD VSS scs8hd_fill_2
XANTENNA__529__A2N _525_/Y VSS VDD scs8hd_diode_2
XFILLER_0_109 VSS VDD scs8hd_fill_1
XANTENNA__393__A _389_/A VSS VDD scs8hd_diode_2
XANTENNA__529__B1 _527_/X VSS VDD scs8hd_diode_2
XANTENNA__568__A _676_/Q VSS VDD scs8hd_diode_2
X_684_ _681_/CLK _684_/D _684_/Q _365_/X VSS VDD scs8hd_dfrtp_4
XFILLER_18_60 VSS VDD scs8hd_decap_6
XFILLER_18_93 VSS VDD scs8hd_decap_4
XFILLER_38_102 VDD VSS scs8hd_fill_2
XFILLER_22_3 VDD VSS scs8hd_fill_2
XFILLER_39_59 VDD VSS scs8hd_fill_2
XFILLER_39_37 VDD VSS scs8hd_fill_2
XFILLER_29_168 VDD VSS scs8hd_fill_2
XFILLER_29_135 VSS VDD scs8hd_decap_6
XANTENNA__388__A _402_/A VSS VDD scs8hd_diode_2
XFILLER_4_245 VSS VDD scs8hd_decap_8
XFILLER_4_212 VDD VSS scs8hd_fill_2
X_598_ _597_/X _598_/X VSS VDD scs8hd_buf_1
X_667_ _667_/CLK _550_/X _545_/A _386_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__480__B _480_/B VSS VDD scs8hd_diode_2
XPHY_17 VSS VDD scs8hd_decap_3
XPHY_28 VSS VDD scs8hd_decap_3
XANTENNA__572__A1N _567_/Y VSS VDD scs8hd_diode_2
XFILLER_41_27 VDD VSS scs8hd_fill_2
XPHY_39 VSS VDD scs8hd_decap_3
XFILLER_1_204 VSS VDD scs8hd_decap_4
XFILLER_9_7 VDD VSS scs8hd_fill_2
X_383_ _386_/A _383_/X VSS VDD scs8hd_buf_1
X_521_ _516_/Y _517_/Y _516_/A _662_/Q _521_/X VSS VDD scs8hd_o22a_4
X_452_ _452_/A _452_/Y VSS VDD scs8hd_inv_8
XANTENNA__581__A _581_/A VSS VDD scs8hd_diode_2
XANTENNA__491__A _490_/X VSS VDD scs8hd_diode_2
XANTENNA__641__D _457_/X VSS VDD scs8hd_diode_2
XFILLER_36_27 VSS VDD scs8hd_decap_4
XFILLER_22_141 VSS VDD scs8hd_fill_1
XANTENNA__576__A _597_/A VSS VDD scs8hd_diode_2
XANTENNA__592__A1 _588_/Y VSS VDD scs8hd_diode_2
XANTENNA__592__B2 _682_/Q VSS VDD scs8hd_diode_2
XFILLER_26_93 VDD VSS scs8hd_fill_2
XFILLER_26_60 VDD VSS scs8hd_fill_2
XFILLER_9_112 VSS VDD scs8hd_decap_8
XFILLER_9_123 VSS VDD scs8hd_decap_8
XFILLER_13_152 VDD VSS scs8hd_fill_2
X_435_ _518_/A x[31] _435_/X VSS VDD scs8hd_and2_4
X_366_ _366_/A _370_/A VSS VDD scs8hd_buf_1
X_504_ _476_/A x[10] _504_/X VSS VDD scs8hd_and2_4
XANTENNA__647__RESETB _410_/X VSS VDD scs8hd_diode_2
XFILLER_9_178 VSS VDD scs8hd_fill_1
XFILLER_13_196 VSS VDD scs8hd_decap_8
XANTENNA__636__D _437_/Y VSS VDD scs8hd_diode_2
XANTENNA__396__A _401_/A VSS VDD scs8hd_diode_2
XFILLER_12_40 VSS VDD scs8hd_decap_3
XFILLER_12_84 VSS VDD scs8hd_decap_4
X_418_ _417_/A _418_/X VSS VDD scs8hd_buf_1
X_349_ _346_/X _347_/X _349_/X VSS VDD scs8hd_xor2_4
XANTENNA__565__B2 _566_/B VSS VDD scs8hd_diode_2
XFILLER_5_181 VDD VSS scs8hd_fill_2
XPHY_209 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__556__B2 _553_/A VSS VDD scs8hd_diode_2
XANTENNA__556__A1 _552_/Y VSS VDD scs8hd_diode_2
XFILLER_24_225 VDD VSS scs8hd_fill_2
XANTENNA__492__B1 _488_/A VSS VDD scs8hd_diode_2
XFILLER_3_118 VSS VDD scs8hd_decap_4
XFILLER_30_206 VSS VDD scs8hd_decap_4
XFILLER_23_72 VDD VSS scs8hd_fill_2
XFILLER_23_50 VDD VSS scs8hd_fill_2
XFILLER_15_236 VDD VSS scs8hd_fill_2
XANTENNA__573__B _573_/B VSS VDD scs8hd_diode_2
XANTENNA__600__A2N _596_/Y VSS VDD scs8hd_diode_2
XFILLER_2_195 VSS VDD scs8hd_decap_4
XFILLER_2_151 VDD VSS scs8hd_fill_2
XANTENNA__483__B x[7] VSS VDD scs8hd_diode_2
XFILLER_0_32 VDD VSS scs8hd_fill_2
XFILLER_0_98 VSS VDD scs8hd_fill_1
XANTENNA__529__A1N _524_/Y VSS VDD scs8hd_diode_2
XANTENNA__529__B2 _528_/X VSS VDD scs8hd_diode_2
XANTENNA__584__A _583_/X VSS VDD scs8hd_diode_2
X_683_ _681_/CLK _683_/D _683_/Q _367_/X VSS VDD scs8hd_dfrtp_4
XFILLER_34_93 VSS VDD scs8hd_decap_3
XFILLER_34_82 VDD VSS scs8hd_fill_2
XANTENNA__653__CLK _651_/CLK VSS VDD scs8hd_diode_2
XFILLER_38_158 VSS VDD scs8hd_decap_3
XFILLER_38_136 VDD VSS scs8hd_fill_2
XFILLER_15_3 VDD VSS scs8hd_fill_2
XANTENNA__456__B1 _452_/A VSS VDD scs8hd_diode_2
XANTENNA__494__A _491_/X VSS VDD scs8hd_diode_2
XANTENNA__644__D _465_/X VSS VDD scs8hd_diode_2
XANTENNA__695__RESETB _357_/A VSS VDD scs8hd_diode_2
XFILLER_39_49 VSS VDD scs8hd_decap_4
XANTENNA__CTS_buf_1_16_A _CTS_root/X VSS VDD scs8hd_diode_2
XANTENNA__676__CLK _667_/CLK VSS VDD scs8hd_diode_2
XFILLER_35_117 VSS VDD scs8hd_fill_1
XFILLER_29_93 VDD VSS scs8hd_fill_2
XFILLER_29_71 VDD VSS scs8hd_fill_2
XFILLER_29_60 VSS VDD scs8hd_fill_1
X_597_ _597_/A x[23] _597_/X VSS VDD scs8hd_and2_4
X_666_ _667_/CLK _544_/X _666_/Q _387_/X VSS VDD scs8hd_dfrtp_4
XFILLER_28_191 VSS VDD scs8hd_fill_1
XANTENNA__489__A _489_/A VSS VDD scs8hd_diode_2
XFILLER_26_128 VDD VSS scs8hd_fill_2
XANTENNA__639__D _450_/X VSS VDD scs8hd_diode_2
XPHY_18 VSS VDD scs8hd_decap_3
XPHY_29 VSS VDD scs8hd_decap_3
XANTENNA__399__A _401_/A VSS VDD scs8hd_diode_2
X_520_ _519_/X _520_/X VSS VDD scs8hd_buf_1
X_382_ _386_/A _382_/X VSS VDD scs8hd_buf_1
XFILLER_25_172 VSS VDD scs8hd_decap_6
XFILLER_25_161 VSS VDD scs8hd_decap_4
X_451_ _451_/A _449_/X _451_/X VSS VDD scs8hd_xor2_4
XFILLER_15_51 VDD VSS scs8hd_fill_2
XFILLER_15_62 VDD VSS scs8hd_fill_2
XFILLER_17_128 VDD VSS scs8hd_fill_2
XFILLER_31_94 VDD VSS scs8hd_fill_2
XFILLER_31_83 VDD VSS scs8hd_fill_2
X_649_ _651_/CLK _486_/X _649_/Q _407_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__341__A2N _337_/Y VSS VDD scs8hd_diode_2
XANTENNA__643__RESETB _414_/X VSS VDD scs8hd_diode_2
XFILLER_31_175 VSS VDD scs8hd_decap_4
XFILLER_31_164 VSS VDD scs8hd_decap_4
XFILLER_31_120 VDD VSS scs8hd_fill_2
XFILLER_16_172 VDD VSS scs8hd_fill_2
XFILLER_39_231 VDD VSS scs8hd_fill_2
XFILLER_22_131 VDD VSS scs8hd_fill_2
XFILLER_22_186 VSS VDD scs8hd_decap_4
XANTENNA__576__B x[20] VSS VDD scs8hd_diode_2
X_503_ _658_/Q _503_/Y VSS VDD scs8hd_inv_8
XFILLER_42_60 VDD VSS scs8hd_fill_2
XANTENNA__592__A2 _589_/Y VSS VDD scs8hd_diode_2
X_365_ _363_/A _365_/X VSS VDD scs8hd_buf_1
X_434_ _434_/A _434_/B _634_/D VSS VDD scs8hd_xor2_4
XFILLER_9_135 VDD VSS scs8hd_fill_2
XFILLER_9_157 VSS VDD scs8hd_decap_4
XFILLER_13_120 VDD VSS scs8hd_fill_2
XFILLER_3_43 VSS VDD scs8hd_decap_3
XFILLER_36_212 VDD VSS scs8hd_fill_2
XANTENNA__652__D _494_/X VSS VDD scs8hd_diode_2
XFILLER_22_19 VDD VSS scs8hd_fill_2
XFILLER_27_245 VSS VDD scs8hd_decap_8
XFILLER_10_123 VDD VSS scs8hd_fill_2
XFILLER_10_189 VDD VSS scs8hd_fill_2
XANTENNA__587__A _584_/X VSS VDD scs8hd_diode_2
XFILLER_18_212 VDD VSS scs8hd_fill_2
X_348_ _343_/Y _344_/Y _346_/X _347_/X _348_/X VSS VDD scs8hd_a2bb2o_4
X_417_ _417_/A _417_/X VSS VDD scs8hd_buf_1
XANTENNA__497__A _476_/A VSS VDD scs8hd_diode_2
XANTENNA__647__D _479_/X VSS VDD scs8hd_diode_2
XFILLER_17_19 VSS VDD scs8hd_decap_4
XANTENNA__556__A2 _553_/Y VSS VDD scs8hd_diode_2
XFILLER_24_215 VSS VDD scs8hd_decap_3
XANTENNA__492__B2 _489_/A VSS VDD scs8hd_diode_2
XANTENNA__492__A1 _488_/Y VSS VDD scs8hd_diode_2
XFILLER_23_62 VDD VSS scs8hd_fill_2
XFILLER_23_40 VSS VDD scs8hd_decap_3
XANTENNA__600__A1N _595_/Y VSS VDD scs8hd_diode_2
XFILLER_17_7 VSS VDD scs8hd_decap_3
XFILLER_9_31 VSS VDD scs8hd_fill_1
XFILLER_28_18 VDD VSS scs8hd_fill_2
XANTENNA__691__RESETB _356_/X VSS VDD scs8hd_diode_2
XFILLER_20_251 VDD VSS scs8hd_fill_2
X_682_ _681_/CLK _601_/X _682_/Q _368_/X VSS VDD scs8hd_dfrtp_4
XFILLER_18_40 VSS VDD scs8hd_fill_1
XFILLER_18_73 VDD VSS scs8hd_fill_2
XFILLER_7_211 VSS VDD scs8hd_decap_4
XANTENNA__456__B2 _644_/Q VSS VDD scs8hd_diode_2
XANTENNA__456__A1 _452_/Y VSS VDD scs8hd_diode_2
XANTENNA__494__B _492_/X VSS VDD scs8hd_diode_2
XFILLER_38_148 VSS VDD scs8hd_fill_1
XANTENNA__638__RESETB _420_/X VSS VDD scs8hd_diode_2
XANTENNA__660__D _660_/D VSS VDD scs8hd_diode_2
XFILLER_29_115 VSS VDD scs8hd_decap_6
XFILLER_37_181 VDD VSS scs8hd_fill_2
XFILLER_4_225 VDD VSS scs8hd_fill_2
XFILLER_20_63 VDD VSS scs8hd_fill_2
X_665_ _667_/CLK _543_/X _538_/A _389_/X VSS VDD scs8hd_dfrtp_4
XANTENNA__595__A _595_/A VSS VDD scs8hd_diode_2
XFILLER_28_170 VDD VSS scs8hd_fill_2
X_596_ _684_/Q _596_/Y VSS VDD scs8hd_inv_8
XFILLER_6_32 VDD VSS scs8hd_fill_2
XFILLER_34_184 VDD VSS scs8hd_fill_2
XANTENNA__655__D _507_/X VSS VDD scs8hd_diode_2
XPHY_19 VSS VDD scs8hd_decap_3
XFILLER_19_181 VDD VSS scs8hd_fill_2
XFILLER_1_228 VDD VSS scs8hd_fill_2
XFILLER_17_118 VSS VDD scs8hd_decap_4
XFILLER_40_154 VSS VDD scs8hd_decap_4
XFILLER_40_143 VDD VSS scs8hd_fill_2
X_381_ _402_/A _386_/A VSS VDD scs8hd_buf_1
XFILLER_25_184 VDD VSS scs8hd_fill_2
XFILLER_25_140 VSS VDD scs8hd_fill_1
X_450_ _445_/Y _446_/Y _451_/A _449_/X _450_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_15_96 VDD VSS scs8hd_fill_2
XANTENNA__643__CLK _648_/CLK VSS VDD scs8hd_diode_2
XFILLER_31_73 VDD VSS scs8hd_fill_2
XFILLER_31_62 VDD VSS scs8hd_fill_2
XANTENNA__341__A1N _336_/Y VSS VDD scs8hd_diode_2
XFILLER_31_110 VDD VSS scs8hd_fill_2
X_648_ _648_/CLK _480_/X _648_/Q _408_/X VSS VDD scs8hd_dfrtp_4
XFILLER_16_151 VDD VSS scs8hd_fill_2
XPHY_190 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__347__B1 _343_/A VSS VDD scs8hd_diode_2
X_579_ _574_/Y _575_/Y _580_/A _578_/X _579_/X VSS VDD scs8hd_a2bb2o_4
XFILLER_39_243 VSS VDD scs8hd_fill_1
XFILLER_39_210 VSS VDD scs8hd_decap_4
XANTENNA__666__CLK _667_/CLK VSS VDD scs8hd_diode_2
XANTENNA__586__B1 _584_/X VSS VDD scs8hd_diode_2
XFILLER_22_154 VDD VSS scs8hd_fill_2
X_CTS_buf_1_48 _CTS_root/X _681_/CLK VSS VDD scs8hd_clkbuf_4
XFILLER_26_84 VSS VDD scs8hd_decap_4
X_502_ _502_/A _502_/Y VSS VDD scs8hd_inv_8
X_433_ _426_/Y _427_/Y _434_/A _434_/B _633_/D VSS VDD scs8hd_a2bb2o_4
XFILLER_42_94 VDD VSS scs8hd_fill_2
XFILLER_13_165 VSS VDD scs8hd_decap_4
X_364_ _363_/A _364_/X VSS VDD scs8hd_buf_1
XANTENNA__689__CLK _681_/CLK VSS VDD scs8hd_diode_2
XFILLER_27_235 VDD VSS scs8hd_fill_2
XFILLER_27_213 VDD VSS scs8hd_fill_2
XFILLER_42_249 VSS VDD scs8hd_decap_4
XFILLER_42_238 VSS VDD scs8hd_decap_8
XFILLER_5_3 VDD VSS scs8hd_fill_2
XFILLER_12_53 VDD VSS scs8hd_fill_2
XANTENNA__686__RESETB _363_/X VSS VDD scs8hd_diode_2
XANTENNA__587__B _587_/B VSS VDD scs8hd_diode_2
X_416_ _373_/A _417_/A VSS VDD scs8hd_buf_1
X_347_ _343_/Y _344_/Y _343_/A _344_/A _347_/X VSS VDD scs8hd_o22a_4
XFILLER_38_3 VDD VSS scs8hd_fill_2
XFILLER_5_172 VDD VSS scs8hd_fill_2
XANTENNA__497__B x[9] VSS VDD scs8hd_diode_2
XANTENNA__663__D _536_/X VSS VDD scs8hd_diode_2
XANTENNA__492__A2 _489_/Y VSS VDD scs8hd_diode_2
XFILLER_15_249 VSS VDD scs8hd_decap_4
XANTENNA__598__A _597_/X VSS VDD scs8hd_diode_2
XFILLER_0_12 VSS VDD scs8hd_decap_12
XFILLER_0_45 VDD VSS scs8hd_fill_2
XFILLER_0_67 VDD VSS scs8hd_fill_2
XFILLER_9_43 VSS VDD scs8hd_decap_12
XANTENNA__658__D _515_/X VSS VDD scs8hd_diode_2
XANTENNA__634__RESETB _424_/X VSS VDD scs8hd_diode_2
X_681_ _681_/CLK _600_/X _595_/A _369_/X VSS VDD scs8hd_dfrtp_4
XFILLER_7_245 VDD VSS scs8hd_fill_2
XFILLER_38_116 VDD VSS scs8hd_fill_2
XANTENNA__456__A2 _453_/Y VSS VDD scs8hd_diode_2
XFILLER_4_215 VSS VDD scs8hd_decap_3
XFILLER_20_20 VDD VSS scs8hd_fill_2
XFILLER_29_62 VDD VSS scs8hd_fill_2
X_595_ _595_/A _595_/Y VSS VDD scs8hd_inv_8
X_664_ _651_/CLK _537_/X _664_/Q _390_/X VSS VDD scs8hd_dfrtp_4
XFILLER_6_11 VSS VDD scs8hd_decap_3
XFILLER_6_99 VSS VDD scs8hd_decap_12
XANTENNA__565__A2N _560_/Y VSS VDD scs8hd_diode_2
XFILLER_20_3 VDD VSS scs8hd_fill_2
XANTENNA__671__D _565_/X VSS VDD scs8hd_diode_2
XFILLER_40_188 VDD VSS scs8hd_fill_2
XFILLER_40_177 VSS VDD scs8hd_decap_4
X_380_ _375_/A _380_/X VSS VDD scs8hd_buf_1
XFILLER_15_31 VDD VSS scs8hd_fill_2
X_647_ _648_/CLK _479_/X _473_/A _410_/X VSS VDD scs8hd_dfrtp_4
XFILLER_16_163 VSS VDD scs8hd_decap_6
XFILLER_16_196 VSS VDD scs8hd_decap_8
X_578_ _574_/Y _575_/Y _574_/A _678_/Q _578_/X VSS VDD scs8hd_o22a_4
XFILLER_31_155 VDD VSS scs8hd_fill_2
XPHY_191 VSS VDD scs8hd_tapvpwrvgnd_1
XPHY_180 VSS VDD scs8hd_tapvpwrvgnd_1
XANTENNA__347__A1 _343_/Y VSS VDD scs8hd_diode_2
XANTENNA__347__B2 _344_/A VSS VDD scs8hd_diode_2
.ends

